localparam
    kMCA_e_brk0                       = 9'h00,
    kMCA_e_clcsec0                    = 9'h01,
    kMCA_e_map0                       = 9'h02,
    kMCA_e_map1                       = 9'h03,
    kMCA_e_map2                       = 9'h04,
    kMCA_e_map3                       = 9'h05,
    kMCA_e_cli0                       = 9'h06,
    kMCA_e_sei0                       = 9'h07,
    kMCA_e_clv0                       = 9'h08,
    kMCA_e_cldsed0                    = 9'h09,
    kMCA_e_clesee0                    = 9'h0A,
    kMCA_e_fetch0                     = 9'h0B,
    kMCA_e_txa0                       = 9'h0C,
    kMCA_e_tya0                       = 9'h0D,
    kMCA_e_txs0                       = 9'h0E,
    kMCA_e_tay0                       = 9'h0F,
    kMCA_e_tax0                       = 9'h10,
    kMCA_e_tsx0                       = 9'h11,
    kMCA_e_tsy0                       = 9'h12,
    kMCA_e_tys0                       = 9'h13,
    kMCA_e_taz0                       = 9'h14,
    kMCA_e_tza0                       = 9'h15,
    kMCA_e_tab0                       = 9'h16,
    kMCA_e_tba0                       = 9'h17,
    kMCA_e_jmp0                       = 9'h18,
    kMCA_e_jmpind0                    = 9'h19,
    kMCA_e_jmpindx0                   = 9'h1A,
    kMCA_e_bra                        = 9'h1B,
    kMCA_e_bpl0                       = 9'h1C,
    kMCA_e_bpl1                       = 9'h1D,
    kMCA_e_bpl2                       = 9'h1E,
    kMCA_e_bmi0                       = 9'h1F,
    kMCA_e_bmi1                       = 9'h20,
    kMCA_e_bmi2                       = 9'h21,
    kMCA_e_bvc0                       = 9'h22,
    kMCA_e_bvc1                       = 9'h23,
    kMCA_e_bvc2                       = 9'h24,
    kMCA_e_bvs0                       = 9'h25,
    kMCA_e_bvs1                       = 9'h26,
    kMCA_e_bvs2                       = 9'h27,
    kMCA_e_bcc0                       = 9'h28,
    kMCA_e_bcc1                       = 9'h29,
    kMCA_e_bcc2                       = 9'h2A,
    kMCA_e_bcs0                       = 9'h2B,
    kMCA_e_bcs1                       = 9'h2C,
    kMCA_e_bcs2                       = 9'h2D,
    kMCA_e_bne0                       = 9'h2E,
    kMCA_e_bne1                       = 9'h2F,
    kMCA_e_bne2                       = 9'h30,
    kMCA_e_beq0                       = 9'h31,
    kMCA_e_beq1                       = 9'h32,
    kMCA_e_beq2                       = 9'h33,
    kMCA_e_braw0                      = 9'h34,
    kMCA_e_deca                       = 9'h35,
    kMCA_e_decx                       = 9'h36,
    kMCA_e_decy                       = 9'h37,
    kMCA_e_decz                       = 9'h38,
    kMCA_e_inca                       = 9'h39,
    kMCA_e_incx                       = 9'h3A,
    kMCA_e_incy                       = 9'h3B,
    kMCA_e_incz                       = 9'h3C,
    kMCA_e_cmpai                      = 9'h3D,
    kMCA_e_cmpxi                      = 9'h3E,
    kMCA_e_cmpyi                      = 9'h3F,
    kMCA_e_cmpzi                      = 9'h40,
    kMCA_e_ldai                       = 9'h41,
    kMCA_e_ldxi                       = 9'h42,
    kMCA_e_ldyi                       = 9'h43,
    kMCA_e_ldzi                       = 9'h44,
    kMCA_e_adci                       = 9'h45,
    kMCA_e_sbci                       = 9'h46,
    kMCA_e_orai                       = 9'h47,
    kMCA_e_andi                       = 9'h48,
    kMCA_e_eori                       = 9'h49,
    kMCA_e_biti                       = 9'h4A,
    kMCA_e_asl_a                      = 9'h4B,
    kMCA_e_rol_a                      = 9'h4C,
    kMCA_e_lsr_a                      = 9'h4D,
    kMCA_e_ror_a                      = 9'h4E,
    kMCA_e_asr_a                      = 9'h4F,
    kMCA_e_push_p                     = 9'h50,
    kMCA_e_push_a                     = 9'h51,
    kMCA_e_push_x                     = 9'h52,
    kMCA_e_push_y                     = 9'h53,
    kMCA_e_push_z                     = 9'h54,
    kMCA_e_pull0                      = 9'h55,
    kMCA_n_pull0                      = 9'h56,
    kMCA_n_pull1                      = 9'h57,
    kMCA_e_jsr0                       = 9'h58,
    kMCA_n_jsr0                       = 9'h59,
    kMCA_e_bsr0                       = 9'h5A,
    kMCA_e_rts0                       = 9'h5B,
    kMCA_e_rti0                       = 9'h5C,
    kMCA_e_jsrind0                    = 9'h5D,
    kMCA_e_jsrindx0                   = 9'h5E,
    kMCA_e_rtn0                       = 9'h5F,
    kMCA_e_inw0                       = 9'h60,
    kMCA_e_dew0                       = 9'h61,
    kMCA_e_asw0                       = 9'h62,
    kMCA_e_row0                       = 9'h63,
    kMCA_e_phwi0                      = 9'h64,
    kMCA_e_phw0                       = 9'h65,
    kMCA_e_neg                        = 9'h66,
    kMCA_e_addr_r_abs0                = 9'h67,
    kMCA_e_addr_r_absx0               = 9'h68,
    kMCA_e_addr_r_absy0               = 9'h69,
    kMCA_n_addr_r_absx0               = 9'h6A,
    kMCA_n_addr_r_absy0               = 9'h6B,
    kMCA_n_addr_m_absx0               = 9'h6C,
    kMCA_n_addr_m_absy0               = 9'h6D,
    kMCA_e_addr_r_zp0                 = 9'h6E,
    kMCA_e_addr_r_zpx0                = 9'h6F,
    kMCA_e_addr_r_zpy0                = 9'h70,
    kMCA_e_addr_r_zpxind0             = 9'h71,
    kMCA_e_addr_r_zpindy0             = 9'h72,
    kMCA_e_addr_r_zpindz0             = 9'h73,
    kMCA_n_addr_r_zpindy0             = 9'h74,
    kMCA_n_addr_r_zpx0                = 9'h75,
    kMCA_n_addr_r_zpx1                = 9'h76,
    kMCA_n_addr_r_zpy0                = 9'h77,
    kMCA_n_addr_r_zpy1                = 9'h78,
    kMCA_n_addr_m_zp0                 = 9'h79,
    kMCA_n_addr_m_abs0                = 9'h7A,
    kMCA_n_addr_m_abs1                = 9'h7B,
    kMCA_n_addr_r_zpxind0             = 9'h7C,
    kMCA_e_addr_spind0                = 9'h7D,
    kMCA_e_addr_w_abs0                = 9'h7E,
    kMCA_e_addr_w_absx0               = 9'h7F,
    kMCA_e_addr_w_absy0               = 9'h80,
    kMCA_n_addr_w_absx0               = 9'h81,
    kMCA_n_addr_w_absy0               = 9'h82,
    kMCA_e_addr_w_zp0_a               = 9'h83,
    kMCA_e_addr_w_zp0_x               = 9'h84,
    kMCA_e_addr_w_zp0_y               = 9'h85,
    kMCA_e_addr_w_zp0_z               = 9'h86,
    kMCA_e_addr_w_zpx0_a              = 9'h87,
    kMCA_e_addr_w_zpx0_y              = 9'h88,
    kMCA_e_addr_w_zpx0_z              = 9'h89,
    kMCA_e_addr_w_zpy0_x              = 9'h8A,
    kMCA_n_addr_w_zpx0                = 9'h8B,
    kMCA_n_addr_w_zpx1_a              = 9'h8C,
    kMCA_n_addr_w_zpx1_y              = 9'h8D,
    kMCA_n_addr_w_zpy0                = 9'h8E,
    kMCA_n_addr_w_zpy1_x              = 9'h8F,
    kMCA_e_addr_w_zpxind0             = 9'h90,
    kMCA_e_addr_w_zpindy0             = 9'h91,
    kMCA_e_addr_w_zpindz0             = 9'h92,
    kMCA_n_addr_m_zpx0                = 9'h93,
    kMCA_n_addr_m_zpx1                = 9'h94,
    kMCA_n_addr_w_zpxind0             = 9'h95,
    kMCA_n_addr_w_zpindy0             = 9'h96,
    kMCA_e_jmp1                       = 9'h97,
    kMCA_e_jmpind1                    = 9'h98,
    kMCA_e_jmpind2                    = 9'h99,
    kMCA_e_jmpind3                    = 9'h9A,
    kMCA_e_jmpindx1                   = 9'h9B,
    kMCA_e_jmpindx2                   = 9'h9C,
    kMCA_e_jmpindx3                   = 9'h9D,
    kMCA_e_bitm1                      = 9'h9E,
    kMCA_e_mem_fetch                  = 9'h9F,
    kMCA_e_push1                      = 9'hA0,
    kMCA_n_jsr1                       = 9'hA1,
    kMCA_e_jsr1                       = 9'hA2,
    kMCA_e_jsr2                       = 9'hA3,
    kMCA_e_jsr3                       = 9'hA4,
    kMCA_e_rts1                       = 9'hA5,
    kMCA_e_rts2                       = 9'hA6,
    kMCA_e_rti1                       = 9'hA7,
    kMCA_e_rti2                       = 9'hA8,
    kMCA_e_rti3                       = 9'hA9,
    kMCA_e_bsr1                       = 9'hAA,
    kMCA_e_bsr2                       = 9'hAB,
    kMCA_e_bsr3                       = 9'hAC,
    kMCA_e_jsrind1                    = 9'hAD,
    kMCA_e_jsrind2                    = 9'hAE,
    kMCA_e_jsrind3                    = 9'hAF,
    kMCA_e_jsrind4                    = 9'hB0,
    kMCA_e_jsrind5                    = 9'hB1,
    kMCA_e_jsrindx1                   = 9'hB2,
    kMCA_e_jsrindx2                   = 9'hB3,
    kMCA_e_jsrindx3                   = 9'hB4,
    kMCA_e_jsrindx4                   = 9'hB5,
    kMCA_e_jsrindx5                   = 9'hB6,
    kMCA_e_rtn1                       = 9'hB7,
    kMCA_e_rtn2                       = 9'hB8,
    kMCA_e_rtn3                       = 9'hB9,
    kMCA_e_rtn4                       = 9'hBA,
    kMCA_e_rtn5                       = 9'hBB,
    kMCA_e_inw1                       = 9'hBC,
    kMCA_e_inw2                       = 9'hBD,
    kMCA_e_inw3                       = 9'hBE,
    kMCA_e_dew1                       = 9'hBF,
    kMCA_e_dew2                       = 9'hC0,
    kMCA_e_dew3                       = 9'hC1,
    kMCA_e_asw1                       = 9'hC2,
    kMCA_e_asw2                       = 9'hC3,
    kMCA_e_asw3                       = 9'hC4,
    kMCA_e_asw4                       = 9'hC5,
    kMCA_e_row1                       = 9'hC6,
    kMCA_e_row2                       = 9'hC7,
    kMCA_e_row3                       = 9'hC8,
    kMCA_e_row4                       = 9'hC9,
    kMCA_e_phwi1                      = 9'hCA,
    kMCA_e_phwi2                      = 9'hCB,
    kMCA_e_phwi3                      = 9'hCC,
    kMCA_e_phw1                       = 9'hCD,
    kMCA_e_phw2                       = 9'hCE,
    kMCA_e_phw3                       = 9'hCF,
    kMCA_e_phw4                       = 9'hD0,
    kMCA_e_phw5                       = 9'hD1,
    kMCA_e_bbr1                       = 9'hD2,
    kMCA_e_bbr2                       = 9'hD3,
    kMCA_e_bbs1                       = 9'hD4,
    kMCA_e_bbs2                       = 9'hD5,
    kMCA_e_trb1                       = 9'hD6,
    kMCA_e_tsb1                       = 9'hD7,
    kMCA_e_addr_r_abs1                = 9'hD8,
    kMCA_e_addr_r_absx1               = 9'hD9,
    kMCA_e_addr_r_absy1               = 9'hDA,
    kMCA_n_addr_r_absx1               = 9'hDB,
    kMCA_n_addr_r_absx2               = 9'hDC,
    kMCA_n_addr_m_absx1               = 9'hDD,
    kMCA_n_addr_m_absx2               = 9'hDE,
    kMCA_n_addr_r_absy1               = 9'hDF,
    kMCA_n_addr_r_absy2               = 9'hE0,
    kMCA_n_addr_m_absy1               = 9'hE1,
    kMCA_n_addr_m_absy2               = 9'hE2,
    kMCA_e_addr_r_zpxind1             = 9'hE3,
    kMCA_e_addr_r_zpxind2             = 9'hE4,
    kMCA_e_addr_w_zpxind1             = 9'hE5,
    kMCA_e_addr_w_zpxind2             = 9'hE6,
    kMCA_e_addr_r_zpindy1             = 9'hE7,
    kMCA_e_addr_r_zpindy2             = 9'hE8,
    kMCA_e_addr_w_zpindy1             = 9'hE9,
    kMCA_e_addr_w_zpindy2             = 9'hEA,
    kMCA_e_addr_r_zpindz1             = 9'hEB,
    kMCA_e_addr_r_zpindz2             = 9'hEC,
    kMCA_e_addr_w_zpindz1             = 9'hED,
    kMCA_e_addr_w_zpindz2             = 9'hEE,
    kMCA_e_addr_spind1                = 9'hEF,
    kMCA_e_addr_spind2                = 9'hF0,
    kMCA_n_addr_r_zpxind1             = 9'hF1,
    kMCA_n_addr_r_zpxind2             = 9'hF2,
    kMCA_n_addr_r_zpxind3             = 9'hF3,
    kMCA_n_addr_w_zpxind1             = 9'hF4,
    kMCA_n_addr_w_zpxind2             = 9'hF5,
    kMCA_n_addr_w_zpxind3             = 9'hF6,
    kMCA_n_addr_r_zpindy1             = 9'hF7,
    kMCA_n_addr_r_zpindy2             = 9'hF8,
    kMCA_n_addr_r_zpindy3             = 9'hF9,
    kMCA_n_addr_w_zpindy1             = 9'hFA,
    kMCA_n_addr_w_zpindy2             = 9'hFB,
    kMCA_n_addr_w_zpindy3             = 9'hFC,
    kMCA_e_brk1                       = 9'hFD,
    kMCA_e_brk2                       = 9'hFE,
    kMCA_e_brk3                       = 9'hFF,
    kMCA_e_brk4                       = 9'h100,
    kMCA_e_brk5                       = 9'h101,
    kMCA_e_addr_r_spind3              = 9'h102,
    kMCA_e_addr_w_abs1_a              = 9'h103,
    kMCA_e_addr_w_abs1_x              = 9'h104,
    kMCA_e_addr_w_abs1_y              = 9'h105,
    kMCA_e_addr_w_abs1_z              = 9'h106,
    kMCA_e_addr_w_absx1_a             = 9'h107,
    kMCA_e_addr_w_absx1_y             = 9'h108,
    kMCA_e_addr_w_absx1_z             = 9'h109,
    kMCA_e_addr_w_absy1_a             = 9'h10A,
    kMCA_e_addr_w_absy1_x             = 9'h10B,
    kMCA_n_addr_w_absx1               = 9'h10C,
    kMCA_n_addr_w_absy1               = 9'h10D,
    kMCA_n_addr_w_absx2_a             = 9'h10E,
    kMCA_n_addr_w_absx2_y             = 9'h10F,
    kMCA_n_addr_w_absx2_z             = 9'h110,
    kMCA_n_addr_w_absy2_a             = 9'h111,
    kMCA_n_addr_w_absy2_x             = 9'h112,
    kMCA_e_addr_w_spind3              = 9'h113,
    kMCA_e_cmpa                       = 9'h114,
    kMCA_e_cmpx                       = 9'h115,
    kMCA_e_cmpy                       = 9'h116,
    kMCA_e_cmpz                       = 9'h117,
    kMCA_e_lda                        = 9'h118,
    kMCA_e_ldx                        = 9'h119,
    kMCA_e_ldy                        = 9'h11A,
    kMCA_e_ldz                        = 9'h11B,
    kMCA_e_adc                        = 9'h11C,
    kMCA_e_sbc                        = 9'h11D,
    kMCA_e_ora                        = 9'h11E,
    kMCA_e_and                        = 9'h11F,
    kMCA_e_eor                        = 9'h120,
    kMCA_e_bitm0                      = 9'h121,
    kMCA_e_asl_mem0                   = 9'h122,
    kMCA_e_rol_mem0                   = 9'h123,
    kMCA_e_lsr_mem0                   = 9'h124,
    kMCA_e_ror_mem0                   = 9'h125,
    kMCA_e_asr_mem0                   = 9'h126,
    kMCA_n_rmw_mem0                   = 9'h127,
    kMCA_e_pull_p                     = 9'h128,
    kMCA_e_pull_a                     = 9'h129,
    kMCA_e_pull_x                     = 9'h12A,
    kMCA_e_pull_y                     = 9'h12B,
    kMCA_e_pull_z                     = 9'h12C,
    kMCA_e_bbr0                       = 9'h12D,
    kMCA_e_bbs0                       = 9'h12E,
    kMCA_e_trb0                       = 9'h12F,
    kMCA_e_tsb0                       = 9'h130,
    kMCA_e_rmb0                       = 9'h131,
    kMCA_e_smb0                       = 9'h132,
    kMCA_e_bplw1                      = 9'h133,
    kMCA_e_bmiw1                      = 9'h134,
    kMCA_e_bvcw1                      = 9'h135,
    kMCA_e_bvsw1                      = 9'h136,
    kMCA_e_braw1                      = 9'h137,
    kMCA_e_bccw1                      = 9'h138,
    kMCA_e_bcsw1                      = 9'h139,
    kMCA_e_bnew1                      = 9'h13A,
    kMCA_e_beqw1                      = 9'h13B,
    kMCA_e_inc_mem0                   = 9'h13C,
    kMCA_e_dec_mem0                   = 9'h13D,
    kMCA_end                          = 9'h13E;
