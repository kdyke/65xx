module memory(clk, we, addr_r, addr_w, di, do);
input clk;
input we;
input [15:0] addr_r;
input [15:0] addr_w;
input [7:0] di;
output [7:0] do;
reg [7:0] ram [0:65535];reg [7:0] do;

initial
begin
ram[16'h000a] = 8'h00; ram[16'h000b] = 8'h00; ram[16'h000c] = 8'h00; ram[16'h000d] = 8'h00; ram[16'h000e] = 8'h00; ram[16'h000f] = 8'h00; ram[16'h0010] = 8'h00; ram[16'h0011] = 8'h00; 
ram[16'h0012] = 8'h00; ram[16'h0013] = 8'hc3; ram[16'h0014] = 8'h82; ram[16'h0015] = 8'h41; ram[16'h0016] = 8'h00; ram[16'h0017] = 8'h7f; ram[16'h0018] = 8'h00; ram[16'h0019] = 8'h1f; 
ram[16'h001a] = 8'h71; ram[16'h001b] = 8'h80; ram[16'h001c] = 8'h0f; ram[16'h001d] = 8'hff; ram[16'h001e] = 8'h7f; ram[16'h001f] = 8'h80; 
ram[16'h0020] = 8'hff; ram[16'h0021] = 8'h0f; ram[16'h0022] = 8'h8f; ram[16'h0023] = 8'h8f; ram[16'h0024] = 8'h10; ram[16'h0025] = 8'h02; ram[16'h0026] = 8'h11; ram[16'h0027] = 8'h02; 
ram[16'h0028] = 8'h12; ram[16'h0029] = 8'h02; ram[16'h002a] = 8'h13; ram[16'h002b] = 8'h02; ram[16'h002c] = 8'h14; ram[16'h002d] = 8'h02; ram[16'h002e] = 8'h18; ram[16'h002f] = 8'h01; 
ram[16'h0030] = 8'h05; ram[16'h0031] = 8'h02; ram[16'h0032] = 8'h06; ram[16'h0033] = 8'h02; ram[16'h0034] = 8'h07; ram[16'h0035] = 8'h02; ram[16'h0036] = 8'h08; ram[16'h0037] = 8'h02; 
ram[16'h0038] = 8'h0d; ram[16'h0039] = 8'h01; ram[16'h003a] = 8'h47; ram[16'h003b] = 8'h02; ram[16'h003c] = 8'h48; ram[16'h003d] = 8'h02; ram[16'h003e] = 8'h49; ram[16'h003f] = 8'h02; 

ram[16'h0040] = 8'h4a; ram[16'h0041] = 8'h02; ram[16'h0042] = 8'h4b; ram[16'h0043] = 8'h02; ram[16'h0044] = 8'h4c; ram[16'h0045] = 8'h02; ram[16'h0046] = 8'h4d; ram[16'h0047] = 8'h02; 
ram[16'h0048] = 8'h4e; ram[16'h0049] = 8'h02; ram[16'h004a] = 8'h43; ram[16'h004b] = 8'h02; ram[16'h004c] = 8'h44; ram[16'h004d] = 8'h02; ram[16'h004e] = 8'h45; ram[16'h004f] = 8'h02; 
ram[16'h0050] = 8'h46; ram[16'h0051] = 8'h02; ram[16'h0052] = 8'h05; ram[16'h0053] = 8'h02; ram[16'h0054] = 8'h06; ram[16'h0055] = 8'h02; ram[16'h0056] = 8'h06; ram[16'h0057] = 8'h01; 
ram[16'h0058] = 8'h07; ram[16'h0059] = 8'h01; 
ram[16'h0200] = 8'h00; ram[16'h0201] = 8'h00; ram[16'h0202] = 8'h00; ram[16'h0203] = 8'h00; ram[16'h0204] = 8'h00; ram[16'h0205] = 8'h00; ram[16'h0206] = 8'h00; ram[16'h0207] = 8'h00; 
ram[16'h0208] = 8'h00; ram[16'h0209] = 8'h00; ram[16'h020a] = 8'h69; ram[16'h020b] = 8'h00; ram[16'h020c] = 8'h60; ram[16'h020d] = 8'he9; ram[16'h020e] = 8'h00; ram[16'h020f] = 8'h60; 
ram[16'h0210] = 8'hc3; ram[16'h0211] = 8'h82; ram[16'h0212] = 8'h41; ram[16'h0213] = 8'h00; ram[16'h0214] = 8'h7f; ram[16'h0215] = 8'h80; ram[16'h0216] = 8'h80; ram[16'h0217] = 8'h00; 
ram[16'h0218] = 8'h02; ram[16'h0219] = 8'h86; ram[16'h021a] = 8'h04; ram[16'h021b] = 8'h82; ram[16'h021c] = 8'h00; ram[16'h021d] = 8'h87; ram[16'h021e] = 8'h05; ram[16'h021f] = 8'h83; 

ram[16'h0220] = 8'h01; ram[16'h0221] = 8'h61; ram[16'h0222] = 8'h41; ram[16'h0223] = 8'h20; ram[16'h0224] = 8'h00; ram[16'h0225] = 8'he1; ram[16'h0226] = 8'hc1; ram[16'h0227] = 8'ha0; 
ram[16'h0228] = 8'h80; ram[16'h0229] = 8'h81; ram[16'h022a] = 8'h01; ram[16'h022b] = 8'h80; ram[16'h022c] = 8'h02; ram[16'h022d] = 8'h81; ram[16'h022e] = 8'h01; ram[16'h022f] = 8'h80; 
ram[16'h0230] = 8'h00; ram[16'h0231] = 8'h01; ram[16'h0232] = 8'h00; ram[16'h0233] = 8'h01; ram[16'h0234] = 8'h02; ram[16'h0235] = 8'h81; ram[16'h0236] = 8'h80; ram[16'h0237] = 8'h81; 
ram[16'h0238] = 8'h80; ram[16'h0239] = 8'h7f; ram[16'h023a] = 8'h80; ram[16'h023b] = 8'hff; ram[16'h023c] = 8'h00; ram[16'h023d] = 8'h01; ram[16'h023e] = 8'h00; ram[16'h023f] = 8'h80; 

ram[16'h0240] = 8'h80; ram[16'h0241] = 8'h02; ram[16'h0242] = 8'h00; ram[16'h0243] = 8'h00; ram[16'h0244] = 8'h1f; ram[16'h0245] = 8'h71; ram[16'h0246] = 8'h80; ram[16'h0247] = 8'h0f; 
ram[16'h0248] = 8'hff; ram[16'h0249] = 8'h7f; ram[16'h024a] = 8'h80; ram[16'h024b] = 8'hff; ram[16'h024c] = 8'h0f; ram[16'h024d] = 8'h8f; ram[16'h024e] = 8'h8f; ram[16'h024f] = 8'h00; 
ram[16'h0250] = 8'hf1; ram[16'h0251] = 8'h1f; ram[16'h0252] = 8'h00; ram[16'h0253] = 8'hf0; ram[16'h0254] = 8'hff; ram[16'h0255] = 8'hff; ram[16'h0256] = 8'hff; ram[16'h0257] = 8'hff; 
ram[16'h0258] = 8'hf0; ram[16'h0259] = 8'hf0; ram[16'h025a] = 8'h0f; ram[16'h025b] = 8'h00; ram[16'h025c] = 8'hff; ram[16'h025d] = 8'h7f; ram[16'h025e] = 8'h80; ram[16'h025f] = 8'h02; 

ram[16'h0260] = 8'h80; ram[16'h0261] = 8'h00; ram[16'h0262] = 8'h80; 
ram[16'h0400] = 8'hd8; ram[16'h0401] = 8'ha2; ram[16'h0402] = 8'hff; ram[16'h0403] = 8'h9a; ram[16'h0404] = 8'ha9; ram[16'h0405] = 8'h00; ram[16'h0406] = 8'h8d; ram[16'h0407] = 8'h02; 
ram[16'h0408] = 8'h02; ram[16'h0409] = 8'had; ram[16'h040a] = 8'h02; ram[16'h040b] = 8'h02; ram[16'h040c] = 8'hc9; ram[16'h040d] = 8'h00; ram[16'h040e] = 8'hd0; ram[16'h040f] = 8'hfe; 
ram[16'h0410] = 8'ha9; ram[16'h0411] = 8'h01; ram[16'h0412] = 8'h8d; ram[16'h0413] = 8'h02; ram[16'h0414] = 8'h02; ram[16'h0415] = 8'ha9; ram[16'h0416] = 8'h99; ram[16'h0417] = 8'ha2; 
ram[16'h0418] = 8'hff; ram[16'h0419] = 8'h9a; ram[16'h041a] = 8'ha2; ram[16'h041b] = 8'h55; ram[16'h041c] = 8'hda; ram[16'h041d] = 8'ha2; ram[16'h041e] = 8'haa; ram[16'h041f] = 8'hda; 

ram[16'h0420] = 8'hec; ram[16'h0421] = 8'hfe; ram[16'h0422] = 8'h01; ram[16'h0423] = 8'hd0; ram[16'h0424] = 8'hfe; ram[16'h0425] = 8'hba; ram[16'h0426] = 8'he0; ram[16'h0427] = 8'hfd; 
ram[16'h0428] = 8'hd0; ram[16'h0429] = 8'hfe; ram[16'h042a] = 8'h7a; ram[16'h042b] = 8'hc0; ram[16'h042c] = 8'haa; ram[16'h042d] = 8'hd0; ram[16'h042e] = 8'hfe; ram[16'h042f] = 8'h7a; 
ram[16'h0430] = 8'hc0; ram[16'h0431] = 8'h55; ram[16'h0432] = 8'hd0; ram[16'h0433] = 8'hfe; ram[16'h0434] = 8'hcc; ram[16'h0435] = 8'hff; ram[16'h0436] = 8'h01; ram[16'h0437] = 8'hd0; 
ram[16'h0438] = 8'hfe; ram[16'h0439] = 8'hba; ram[16'h043a] = 8'he0; ram[16'h043b] = 8'hff; ram[16'h043c] = 8'hd0; ram[16'h043d] = 8'hfe; ram[16'h043e] = 8'ha0; ram[16'h043f] = 8'ha5; 

ram[16'h0440] = 8'h5a; ram[16'h0441] = 8'ha0; ram[16'h0442] = 8'h5a; ram[16'h0443] = 8'h5a; ram[16'h0444] = 8'hcc; ram[16'h0445] = 8'hfe; ram[16'h0446] = 8'h01; ram[16'h0447] = 8'hd0; 
ram[16'h0448] = 8'hfe; ram[16'h0449] = 8'hba; ram[16'h044a] = 8'he0; ram[16'h044b] = 8'hfd; ram[16'h044c] = 8'hd0; ram[16'h044d] = 8'hfe; ram[16'h044e] = 8'hfa; ram[16'h044f] = 8'he0; 
ram[16'h0450] = 8'h5a; ram[16'h0451] = 8'hd0; ram[16'h0452] = 8'hfe; ram[16'h0453] = 8'hfa; ram[16'h0454] = 8'he0; ram[16'h0455] = 8'ha5; ram[16'h0456] = 8'hd0; ram[16'h0457] = 8'hfe; 
ram[16'h0458] = 8'hec; ram[16'h0459] = 8'hff; ram[16'h045a] = 8'h01; ram[16'h045b] = 8'hd0; ram[16'h045c] = 8'hfe; ram[16'h045d] = 8'hba; ram[16'h045e] = 8'he0; ram[16'h045f] = 8'hff; 

ram[16'h0460] = 8'hd0; ram[16'h0461] = 8'hfe; ram[16'h0462] = 8'hc9; ram[16'h0463] = 8'h99; ram[16'h0464] = 8'hd0; ram[16'h0465] = 8'hfe; ram[16'h0466] = 8'had; ram[16'h0467] = 8'h02; 
ram[16'h0468] = 8'h02; ram[16'h0469] = 8'hc9; ram[16'h046a] = 8'h01; ram[16'h046b] = 8'hd0; ram[16'h046c] = 8'hfe; ram[16'h046d] = 8'ha9; ram[16'h046e] = 8'h02; ram[16'h046f] = 8'h8d; 
ram[16'h0470] = 8'h02; ram[16'h0471] = 8'h02; ram[16'h0472] = 8'ha0; ram[16'h0473] = 8'haa; ram[16'h0474] = 8'ha9; ram[16'h0475] = 8'hff; ram[16'h0476] = 8'h48; ram[16'h0477] = 8'ha2; 
ram[16'h0478] = 8'h01; ram[16'h0479] = 8'h28; ram[16'h047a] = 8'hda; ram[16'h047b] = 8'h08; ram[16'h047c] = 8'he0; ram[16'h047d] = 8'h01; ram[16'h047e] = 8'hd0; ram[16'h047f] = 8'hfe; 

ram[16'h0480] = 8'h68; ram[16'h0481] = 8'h48; ram[16'h0482] = 8'hc9; ram[16'h0483] = 8'hff; ram[16'h0484] = 8'hd0; ram[16'h0485] = 8'hfe; ram[16'h0486] = 8'h28; ram[16'h0487] = 8'ha9; 
ram[16'h0488] = 8'h00; ram[16'h0489] = 8'h48; ram[16'h048a] = 8'ha2; ram[16'h048b] = 8'h00; ram[16'h048c] = 8'h28; ram[16'h048d] = 8'hda; ram[16'h048e] = 8'h08; ram[16'h048f] = 8'he0; 
ram[16'h0490] = 8'h00; ram[16'h0491] = 8'hd0; ram[16'h0492] = 8'hfe; ram[16'h0493] = 8'h68; ram[16'h0494] = 8'h48; ram[16'h0495] = 8'hc9; ram[16'h0496] = 8'h30; ram[16'h0497] = 8'hd0; 
ram[16'h0498] = 8'hfe; ram[16'h0499] = 8'h28; ram[16'h049a] = 8'ha9; ram[16'h049b] = 8'hff; ram[16'h049c] = 8'h48; ram[16'h049d] = 8'ha2; ram[16'h049e] = 8'hff; ram[16'h049f] = 8'h28; 

ram[16'h04a0] = 8'hda; ram[16'h04a1] = 8'h08; ram[16'h04a2] = 8'he0; ram[16'h04a3] = 8'hff; ram[16'h04a4] = 8'hd0; ram[16'h04a5] = 8'hfe; ram[16'h04a6] = 8'h68; ram[16'h04a7] = 8'h48; 
ram[16'h04a8] = 8'hc9; ram[16'h04a9] = 8'hff; ram[16'h04aa] = 8'hd0; ram[16'h04ab] = 8'hfe; ram[16'h04ac] = 8'h28; ram[16'h04ad] = 8'ha9; ram[16'h04ae] = 8'h00; ram[16'h04af] = 8'h48; 
ram[16'h04b0] = 8'ha2; ram[16'h04b1] = 8'h01; ram[16'h04b2] = 8'h28; ram[16'h04b3] = 8'hda; ram[16'h04b4] = 8'h08; ram[16'h04b5] = 8'he0; ram[16'h04b6] = 8'h01; ram[16'h04b7] = 8'hd0; 
ram[16'h04b8] = 8'hfe; ram[16'h04b9] = 8'h68; ram[16'h04ba] = 8'h48; ram[16'h04bb] = 8'hc9; ram[16'h04bc] = 8'h30; ram[16'h04bd] = 8'hd0; ram[16'h04be] = 8'hfe; ram[16'h04bf] = 8'h28; 

ram[16'h04c0] = 8'ha9; ram[16'h04c1] = 8'hff; ram[16'h04c2] = 8'h48; ram[16'h04c3] = 8'ha2; ram[16'h04c4] = 8'h00; ram[16'h04c5] = 8'h28; ram[16'h04c6] = 8'hda; ram[16'h04c7] = 8'h08; 
ram[16'h04c8] = 8'he0; ram[16'h04c9] = 8'h00; ram[16'h04ca] = 8'hd0; ram[16'h04cb] = 8'hfe; ram[16'h04cc] = 8'h68; ram[16'h04cd] = 8'h48; ram[16'h04ce] = 8'hc9; ram[16'h04cf] = 8'hff; 
ram[16'h04d0] = 8'hd0; ram[16'h04d1] = 8'hfe; ram[16'h04d2] = 8'h28; ram[16'h04d3] = 8'ha9; ram[16'h04d4] = 8'h00; ram[16'h04d5] = 8'h48; ram[16'h04d6] = 8'ha2; ram[16'h04d7] = 8'hff; 
ram[16'h04d8] = 8'h28; ram[16'h04d9] = 8'hda; ram[16'h04da] = 8'h08; ram[16'h04db] = 8'he0; ram[16'h04dc] = 8'hff; ram[16'h04dd] = 8'hd0; ram[16'h04de] = 8'hfe; ram[16'h04df] = 8'h68; 

ram[16'h04e0] = 8'h48; ram[16'h04e1] = 8'hc9; ram[16'h04e2] = 8'h30; ram[16'h04e3] = 8'hd0; ram[16'h04e4] = 8'hfe; ram[16'h04e5] = 8'h28; ram[16'h04e6] = 8'ha9; ram[16'h04e7] = 8'hff; 
ram[16'h04e8] = 8'h48; ram[16'h04e9] = 8'ha2; ram[16'h04ea] = 8'h00; ram[16'h04eb] = 8'h28; ram[16'h04ec] = 8'hfa; ram[16'h04ed] = 8'h08; ram[16'h04ee] = 8'he0; ram[16'h04ef] = 8'hff; 
ram[16'h04f0] = 8'hd0; ram[16'h04f1] = 8'hfe; ram[16'h04f2] = 8'h68; ram[16'h04f3] = 8'h48; ram[16'h04f4] = 8'hc9; ram[16'h04f5] = 8'hfd; ram[16'h04f6] = 8'hd0; ram[16'h04f7] = 8'hfe; 
ram[16'h04f8] = 8'h28; ram[16'h04f9] = 8'ha9; ram[16'h04fa] = 8'h00; ram[16'h04fb] = 8'h48; ram[16'h04fc] = 8'ha2; ram[16'h04fd] = 8'hff; ram[16'h04fe] = 8'h28; ram[16'h04ff] = 8'hfa; 

ram[16'h0500] = 8'h08; ram[16'h0501] = 8'he0; ram[16'h0502] = 8'h00; ram[16'h0503] = 8'hd0; ram[16'h0504] = 8'hfe; ram[16'h0505] = 8'h68; ram[16'h0506] = 8'h48; ram[16'h0507] = 8'hc9; 
ram[16'h0508] = 8'h32; ram[16'h0509] = 8'hd0; ram[16'h050a] = 8'hfe; ram[16'h050b] = 8'h28; ram[16'h050c] = 8'ha9; ram[16'h050d] = 8'hff; ram[16'h050e] = 8'h48; ram[16'h050f] = 8'ha2; 
ram[16'h0510] = 8'hfe; ram[16'h0511] = 8'h28; ram[16'h0512] = 8'hfa; ram[16'h0513] = 8'h08; ram[16'h0514] = 8'he0; ram[16'h0515] = 8'h01; ram[16'h0516] = 8'hd0; ram[16'h0517] = 8'hfe; 
ram[16'h0518] = 8'h68; ram[16'h0519] = 8'h48; ram[16'h051a] = 8'hc9; ram[16'h051b] = 8'h7d; ram[16'h051c] = 8'hd0; ram[16'h051d] = 8'hfe; ram[16'h051e] = 8'h28; ram[16'h051f] = 8'ha9; 

ram[16'h0520] = 8'h00; ram[16'h0521] = 8'h48; ram[16'h0522] = 8'ha2; ram[16'h0523] = 8'h00; ram[16'h0524] = 8'h28; ram[16'h0525] = 8'hfa; ram[16'h0526] = 8'h08; ram[16'h0527] = 8'he0; 
ram[16'h0528] = 8'hff; ram[16'h0529] = 8'hd0; ram[16'h052a] = 8'hfe; ram[16'h052b] = 8'h68; ram[16'h052c] = 8'h48; ram[16'h052d] = 8'hc9; ram[16'h052e] = 8'hb0; ram[16'h052f] = 8'hd0; 
ram[16'h0530] = 8'hfe; ram[16'h0531] = 8'h28; ram[16'h0532] = 8'ha9; ram[16'h0533] = 8'hff; ram[16'h0534] = 8'h48; ram[16'h0535] = 8'ha2; ram[16'h0536] = 8'hff; ram[16'h0537] = 8'h28; 
ram[16'h0538] = 8'hfa; ram[16'h0539] = 8'h08; ram[16'h053a] = 8'he0; ram[16'h053b] = 8'h00; ram[16'h053c] = 8'hd0; ram[16'h053d] = 8'hfe; ram[16'h053e] = 8'h68; ram[16'h053f] = 8'h48; 

ram[16'h0540] = 8'hc9; ram[16'h0541] = 8'h7f; ram[16'h0542] = 8'hd0; ram[16'h0543] = 8'hfe; ram[16'h0544] = 8'h28; ram[16'h0545] = 8'ha9; ram[16'h0546] = 8'h00; ram[16'h0547] = 8'h48; 
ram[16'h0548] = 8'ha2; ram[16'h0549] = 8'hfe; ram[16'h054a] = 8'h28; ram[16'h054b] = 8'hfa; ram[16'h054c] = 8'h08; ram[16'h054d] = 8'he0; ram[16'h054e] = 8'h01; ram[16'h054f] = 8'hd0; 
ram[16'h0550] = 8'hfe; ram[16'h0551] = 8'h68; ram[16'h0552] = 8'h48; ram[16'h0553] = 8'hc9; ram[16'h0554] = 8'h30; ram[16'h0555] = 8'hd0; ram[16'h0556] = 8'hfe; ram[16'h0557] = 8'h28; 
ram[16'h0558] = 8'hc0; ram[16'h0559] = 8'haa; ram[16'h055a] = 8'hd0; ram[16'h055b] = 8'hfe; ram[16'h055c] = 8'had; ram[16'h055d] = 8'h02; ram[16'h055e] = 8'h02; ram[16'h055f] = 8'hc9; 

ram[16'h0560] = 8'h02; ram[16'h0561] = 8'hd0; ram[16'h0562] = 8'hfe; ram[16'h0563] = 8'ha9; ram[16'h0564] = 8'h03; ram[16'h0565] = 8'h8d; ram[16'h0566] = 8'h02; ram[16'h0567] = 8'h02; 
ram[16'h0568] = 8'ha2; ram[16'h0569] = 8'h55; ram[16'h056a] = 8'ha9; ram[16'h056b] = 8'hff; ram[16'h056c] = 8'h48; ram[16'h056d] = 8'ha0; ram[16'h056e] = 8'h01; ram[16'h056f] = 8'h28; 
ram[16'h0570] = 8'h5a; ram[16'h0571] = 8'h08; ram[16'h0572] = 8'hc0; ram[16'h0573] = 8'h01; ram[16'h0574] = 8'hd0; ram[16'h0575] = 8'hfe; ram[16'h0576] = 8'h68; ram[16'h0577] = 8'h48; 
ram[16'h0578] = 8'hc9; ram[16'h0579] = 8'hff; ram[16'h057a] = 8'hd0; ram[16'h057b] = 8'hfe; ram[16'h057c] = 8'h28; ram[16'h057d] = 8'ha9; ram[16'h057e] = 8'h00; ram[16'h057f] = 8'h48; 

ram[16'h0580] = 8'ha0; ram[16'h0581] = 8'h00; ram[16'h0582] = 8'h28; ram[16'h0583] = 8'h5a; ram[16'h0584] = 8'h08; ram[16'h0585] = 8'hc0; ram[16'h0586] = 8'h00; ram[16'h0587] = 8'hd0; 
ram[16'h0588] = 8'hfe; ram[16'h0589] = 8'h68; ram[16'h058a] = 8'h48; ram[16'h058b] = 8'hc9; ram[16'h058c] = 8'h30; ram[16'h058d] = 8'hd0; ram[16'h058e] = 8'hfe; ram[16'h058f] = 8'h28; 
ram[16'h0590] = 8'ha9; ram[16'h0591] = 8'hff; ram[16'h0592] = 8'h48; ram[16'h0593] = 8'ha0; ram[16'h0594] = 8'hff; ram[16'h0595] = 8'h28; ram[16'h0596] = 8'h5a; ram[16'h0597] = 8'h08; 
ram[16'h0598] = 8'hc0; ram[16'h0599] = 8'hff; ram[16'h059a] = 8'hd0; ram[16'h059b] = 8'hfe; ram[16'h059c] = 8'h68; ram[16'h059d] = 8'h48; ram[16'h059e] = 8'hc9; ram[16'h059f] = 8'hff; 

ram[16'h05a0] = 8'hd0; ram[16'h05a1] = 8'hfe; ram[16'h05a2] = 8'h28; ram[16'h05a3] = 8'ha9; ram[16'h05a4] = 8'h00; ram[16'h05a5] = 8'h48; ram[16'h05a6] = 8'ha0; ram[16'h05a7] = 8'h01; 
ram[16'h05a8] = 8'h28; ram[16'h05a9] = 8'h5a; ram[16'h05aa] = 8'h08; ram[16'h05ab] = 8'hc0; ram[16'h05ac] = 8'h01; ram[16'h05ad] = 8'hd0; ram[16'h05ae] = 8'hfe; ram[16'h05af] = 8'h68; 
ram[16'h05b0] = 8'h48; ram[16'h05b1] = 8'hc9; ram[16'h05b2] = 8'h30; ram[16'h05b3] = 8'hd0; ram[16'h05b4] = 8'hfe; ram[16'h05b5] = 8'h28; ram[16'h05b6] = 8'ha9; ram[16'h05b7] = 8'hff; 
ram[16'h05b8] = 8'h48; ram[16'h05b9] = 8'ha0; ram[16'h05ba] = 8'h00; ram[16'h05bb] = 8'h28; ram[16'h05bc] = 8'h5a; ram[16'h05bd] = 8'h08; ram[16'h05be] = 8'hc0; ram[16'h05bf] = 8'h00; 

ram[16'h05c0] = 8'hd0; ram[16'h05c1] = 8'hfe; ram[16'h05c2] = 8'h68; ram[16'h05c3] = 8'h48; ram[16'h05c4] = 8'hc9; ram[16'h05c5] = 8'hff; ram[16'h05c6] = 8'hd0; ram[16'h05c7] = 8'hfe; 
ram[16'h05c8] = 8'h28; ram[16'h05c9] = 8'ha9; ram[16'h05ca] = 8'h00; ram[16'h05cb] = 8'h48; ram[16'h05cc] = 8'ha0; ram[16'h05cd] = 8'hff; ram[16'h05ce] = 8'h28; ram[16'h05cf] = 8'h5a; 
ram[16'h05d0] = 8'h08; ram[16'h05d1] = 8'hc0; ram[16'h05d2] = 8'hff; ram[16'h05d3] = 8'hd0; ram[16'h05d4] = 8'hfe; ram[16'h05d5] = 8'h68; ram[16'h05d6] = 8'h48; ram[16'h05d7] = 8'hc9; 
ram[16'h05d8] = 8'h30; ram[16'h05d9] = 8'hd0; ram[16'h05da] = 8'hfe; ram[16'h05db] = 8'h28; ram[16'h05dc] = 8'ha9; ram[16'h05dd] = 8'hff; ram[16'h05de] = 8'h48; ram[16'h05df] = 8'ha0; 

ram[16'h05e0] = 8'h00; ram[16'h05e1] = 8'h28; ram[16'h05e2] = 8'h7a; ram[16'h05e3] = 8'h08; ram[16'h05e4] = 8'hc0; ram[16'h05e5] = 8'hff; ram[16'h05e6] = 8'hd0; ram[16'h05e7] = 8'hfe; 
ram[16'h05e8] = 8'h68; ram[16'h05e9] = 8'h48; ram[16'h05ea] = 8'hc9; ram[16'h05eb] = 8'hfd; ram[16'h05ec] = 8'hd0; ram[16'h05ed] = 8'hfe; ram[16'h05ee] = 8'h28; ram[16'h05ef] = 8'ha9; 
ram[16'h05f0] = 8'h00; ram[16'h05f1] = 8'h48; ram[16'h05f2] = 8'ha0; ram[16'h05f3] = 8'hff; ram[16'h05f4] = 8'h28; ram[16'h05f5] = 8'h7a; ram[16'h05f6] = 8'h08; ram[16'h05f7] = 8'hc0; 
ram[16'h05f8] = 8'h00; ram[16'h05f9] = 8'hd0; ram[16'h05fa] = 8'hfe; ram[16'h05fb] = 8'h68; ram[16'h05fc] = 8'h48; ram[16'h05fd] = 8'hc9; ram[16'h05fe] = 8'h32; ram[16'h05ff] = 8'hd0; 

ram[16'h0600] = 8'hfe; ram[16'h0601] = 8'h28; ram[16'h0602] = 8'ha9; ram[16'h0603] = 8'hff; ram[16'h0604] = 8'h48; ram[16'h0605] = 8'ha0; ram[16'h0606] = 8'hfe; ram[16'h0607] = 8'h28; 
ram[16'h0608] = 8'h7a; ram[16'h0609] = 8'h08; ram[16'h060a] = 8'hc0; ram[16'h060b] = 8'h01; ram[16'h060c] = 8'hd0; ram[16'h060d] = 8'hfe; ram[16'h060e] = 8'h68; ram[16'h060f] = 8'h48; 
ram[16'h0610] = 8'hc9; ram[16'h0611] = 8'h7d; ram[16'h0612] = 8'hd0; ram[16'h0613] = 8'hfe; ram[16'h0614] = 8'h28; ram[16'h0615] = 8'ha9; ram[16'h0616] = 8'h00; ram[16'h0617] = 8'h48; 
ram[16'h0618] = 8'ha0; ram[16'h0619] = 8'h00; ram[16'h061a] = 8'h28; ram[16'h061b] = 8'h7a; ram[16'h061c] = 8'h08; ram[16'h061d] = 8'hc0; ram[16'h061e] = 8'hff; ram[16'h061f] = 8'hd0; 

ram[16'h0620] = 8'hfe; ram[16'h0621] = 8'h68; ram[16'h0622] = 8'h48; ram[16'h0623] = 8'hc9; ram[16'h0624] = 8'hb0; ram[16'h0625] = 8'hd0; ram[16'h0626] = 8'hfe; ram[16'h0627] = 8'h28; 
ram[16'h0628] = 8'ha9; ram[16'h0629] = 8'hff; ram[16'h062a] = 8'h48; ram[16'h062b] = 8'ha0; ram[16'h062c] = 8'hff; ram[16'h062d] = 8'h28; ram[16'h062e] = 8'h7a; ram[16'h062f] = 8'h08; 
ram[16'h0630] = 8'hc0; ram[16'h0631] = 8'h00; ram[16'h0632] = 8'hd0; ram[16'h0633] = 8'hfe; ram[16'h0634] = 8'h68; ram[16'h0635] = 8'h48; ram[16'h0636] = 8'hc9; ram[16'h0637] = 8'h7f; 
ram[16'h0638] = 8'hd0; ram[16'h0639] = 8'hfe; ram[16'h063a] = 8'h28; ram[16'h063b] = 8'ha9; ram[16'h063c] = 8'h00; ram[16'h063d] = 8'h48; ram[16'h063e] = 8'ha0; ram[16'h063f] = 8'hfe; 

ram[16'h0640] = 8'h28; ram[16'h0641] = 8'h7a; ram[16'h0642] = 8'h08; ram[16'h0643] = 8'hc0; ram[16'h0644] = 8'h01; ram[16'h0645] = 8'hd0; ram[16'h0646] = 8'hfe; ram[16'h0647] = 8'h68; 
ram[16'h0648] = 8'h48; ram[16'h0649] = 8'hc9; ram[16'h064a] = 8'h30; ram[16'h064b] = 8'hd0; ram[16'h064c] = 8'hfe; ram[16'h064d] = 8'h28; ram[16'h064e] = 8'he0; ram[16'h064f] = 8'h55; 
ram[16'h0650] = 8'hd0; ram[16'h0651] = 8'hfe; ram[16'h0652] = 8'had; ram[16'h0653] = 8'h02; ram[16'h0654] = 8'h02; ram[16'h0655] = 8'hc9; ram[16'h0656] = 8'h03; ram[16'h0657] = 8'hd0; 
ram[16'h0658] = 8'hfe; ram[16'h0659] = 8'ha9; ram[16'h065a] = 8'h04; ram[16'h065b] = 8'h8d; ram[16'h065c] = 8'h02; ram[16'h065d] = 8'h02; ram[16'h065e] = 8'ha2; ram[16'h065f] = 8'h81; 

ram[16'h0660] = 8'ha0; ram[16'h0661] = 8'h7e; ram[16'h0662] = 8'ha9; ram[16'h0663] = 8'hff; ram[16'h0664] = 8'h48; ram[16'h0665] = 8'ha9; ram[16'h0666] = 8'h00; ram[16'h0667] = 8'h28; 
ram[16'h0668] = 8'h80; ram[16'h0669] = 8'h03; ram[16'h066a] = 8'h4c; ram[16'h066b] = 8'h6a; ram[16'h066c] = 8'h06; ram[16'h066d] = 8'h08; ram[16'h066e] = 8'hc9; ram[16'h066f] = 8'h00; 
ram[16'h0670] = 8'hd0; ram[16'h0671] = 8'hfe; ram[16'h0672] = 8'h68; ram[16'h0673] = 8'h48; ram[16'h0674] = 8'hc9; ram[16'h0675] = 8'hff; ram[16'h0676] = 8'hd0; ram[16'h0677] = 8'hfe; 
ram[16'h0678] = 8'h28; ram[16'h0679] = 8'ha9; ram[16'h067a] = 8'h00; ram[16'h067b] = 8'h48; ram[16'h067c] = 8'ha9; ram[16'h067d] = 8'hff; ram[16'h067e] = 8'h28; ram[16'h067f] = 8'h80; 

ram[16'h0680] = 8'h03; ram[16'h0681] = 8'h4c; ram[16'h0682] = 8'h81; ram[16'h0683] = 8'h06; ram[16'h0684] = 8'h08; ram[16'h0685] = 8'hc9; ram[16'h0686] = 8'hff; ram[16'h0687] = 8'hd0; 
ram[16'h0688] = 8'hfe; ram[16'h0689] = 8'h68; ram[16'h068a] = 8'h48; ram[16'h068b] = 8'hc9; ram[16'h068c] = 8'h30; ram[16'h068d] = 8'hd0; ram[16'h068e] = 8'hfe; ram[16'h068f] = 8'h28; 
ram[16'h0690] = 8'he0; ram[16'h0691] = 8'h81; ram[16'h0692] = 8'hd0; ram[16'h0693] = 8'hfe; ram[16'h0694] = 8'hc0; ram[16'h0695] = 8'h7e; ram[16'h0696] = 8'hd0; ram[16'h0697] = 8'hfe; 
ram[16'h0698] = 8'had; ram[16'h0699] = 8'h02; ram[16'h069a] = 8'h02; ram[16'h069b] = 8'hc9; ram[16'h069c] = 8'h04; ram[16'h069d] = 8'hd0; ram[16'h069e] = 8'hfe; ram[16'h069f] = 8'ha9; 

ram[16'h06a0] = 8'h05; ram[16'h06a1] = 8'h8d; ram[16'h06a2] = 8'h02; ram[16'h06a3] = 8'h02; ram[16'h06a4] = 8'ha0; ram[16'h06a5] = 8'h00; ram[16'h06a6] = 8'h80; ram[16'h06a7] = 8'h61; 
ram[16'h06a8] = 8'hc0; ram[16'h06a9] = 8'h01; ram[16'h06aa] = 8'hd0; ram[16'h06ab] = 8'hfe; ram[16'h06ac] = 8'hc8; ram[16'h06ad] = 8'h80; ram[16'h06ae] = 8'h53; ram[16'h06af] = 8'hc0; 
ram[16'h06b0] = 8'h03; ram[16'h06b1] = 8'hd0; ram[16'h06b2] = 8'hfe; ram[16'h06b3] = 8'hc8; ram[16'h06b4] = 8'h80; ram[16'h06b5] = 8'h45; ram[16'h06b6] = 8'hc0; ram[16'h06b7] = 8'h05; 
ram[16'h06b8] = 8'hd0; ram[16'h06b9] = 8'hfe; ram[16'h06ba] = 8'hc8; ram[16'h06bb] = 8'ha0; ram[16'h06bc] = 8'h00; ram[16'h06bd] = 8'h80; ram[16'h06be] = 8'h04; ram[16'h06bf] = 8'hc8; 

ram[16'h06c0] = 8'hc8; ram[16'h06c1] = 8'hc8; ram[16'h06c2] = 8'hc8; ram[16'h06c3] = 8'h80; ram[16'h06c4] = 8'h03; ram[16'h06c5] = 8'hc8; ram[16'h06c6] = 8'hc8; ram[16'h06c7] = 8'hc8; 
ram[16'h06c8] = 8'hc8; ram[16'h06c9] = 8'h80; ram[16'h06ca] = 8'h02; ram[16'h06cb] = 8'hc8; ram[16'h06cc] = 8'hc8; ram[16'h06cd] = 8'hc8; ram[16'h06ce] = 8'hc8; ram[16'h06cf] = 8'h80; 
ram[16'h06d0] = 8'h01; ram[16'h06d1] = 8'hc8; ram[16'h06d2] = 8'hc8; ram[16'h06d3] = 8'hc8; ram[16'h06d4] = 8'hc8; ram[16'h06d5] = 8'h80; ram[16'h06d6] = 8'h00; ram[16'h06d7] = 8'hc8; 
ram[16'h06d8] = 8'hc8; ram[16'h06d9] = 8'hc8; ram[16'h06da] = 8'hc8; ram[16'h06db] = 8'hc0; ram[16'h06dc] = 8'h0a; ram[16'h06dd] = 8'hd0; ram[16'h06de] = 8'hfe; ram[16'h06df] = 8'h80; 

ram[16'h06e0] = 8'h12; ram[16'h06e1] = 8'h88; ram[16'h06e2] = 8'h88; ram[16'h06e3] = 8'h88; ram[16'h06e4] = 8'h88; ram[16'h06e5] = 8'h80; ram[16'h06e6] = 8'h0e; ram[16'h06e7] = 8'h88; 
ram[16'h06e8] = 8'h88; ram[16'h06e9] = 8'h88; ram[16'h06ea] = 8'h80; ram[16'h06eb] = 8'hf5; ram[16'h06ec] = 8'h88; ram[16'h06ed] = 8'h88; ram[16'h06ee] = 8'h80; ram[16'h06ef] = 8'hf7; 
ram[16'h06f0] = 8'h88; ram[16'h06f1] = 8'h80; ram[16'h06f2] = 8'hf9; ram[16'h06f3] = 8'h80; ram[16'h06f4] = 8'hfb; ram[16'h06f5] = 8'hc0; ram[16'h06f6] = 8'h00; ram[16'h06f7] = 8'hd0; 
ram[16'h06f8] = 8'hfe; ram[16'h06f9] = 8'h80; ram[16'h06fa] = 8'h15; ram[16'h06fb] = 8'hc0; ram[16'h06fc] = 8'h04; ram[16'h06fd] = 8'hd0; ram[16'h06fe] = 8'hfe; ram[16'h06ff] = 8'hc8; 

ram[16'h0700] = 8'h80; ram[16'h0701] = 8'hb4; ram[16'h0702] = 8'hc0; ram[16'h0703] = 8'h02; ram[16'h0704] = 8'hd0; ram[16'h0705] = 8'hfe; ram[16'h0706] = 8'hc8; ram[16'h0707] = 8'h80; 
ram[16'h0708] = 8'ha6; ram[16'h0709] = 8'hc0; ram[16'h070a] = 8'h00; ram[16'h070b] = 8'hd0; ram[16'h070c] = 8'hfe; ram[16'h070d] = 8'hc8; ram[16'h070e] = 8'h80; ram[16'h070f] = 8'h98; 
ram[16'h0710] = 8'had; ram[16'h0711] = 8'h02; ram[16'h0712] = 8'h02; ram[16'h0713] = 8'hc9; ram[16'h0714] = 8'h05; ram[16'h0715] = 8'hd0; ram[16'h0716] = 8'hfe; ram[16'h0717] = 8'ha9; 
ram[16'h0718] = 8'h06; ram[16'h0719] = 8'h8d; ram[16'h071a] = 8'h02; ram[16'h071b] = 8'h02; ram[16'h071c] = 8'ha2; ram[16'h071d] = 8'h11; ram[16'h071e] = 8'ha0; ram[16'h071f] = 8'h22; 

ram[16'h0720] = 8'ha9; ram[16'h0721] = 8'h01; ram[16'h0722] = 8'h85; ram[16'h0723] = 8'h0c; ram[16'h0724] = 8'ha9; ram[16'h0725] = 8'h00; ram[16'h0726] = 8'h48; ram[16'h0727] = 8'ha9; 
ram[16'h0728] = 8'h33; ram[16'h0729] = 8'h28; ram[16'h072a] = 8'h0f; ram[16'h072b] = 8'h0c; ram[16'h072c] = 8'h06; ram[16'h072d] = 8'h8f; ram[16'h072e] = 8'h0c; ram[16'h072f] = 8'h06; 
ram[16'h0730] = 8'h4c; ram[16'h0731] = 8'h30; ram[16'h0732] = 8'h07; ram[16'h0733] = 8'h4c; ram[16'h0734] = 8'h33; ram[16'h0735] = 8'h07; ram[16'h0736] = 8'h08; ram[16'h0737] = 8'hc9; 
ram[16'h0738] = 8'h33; ram[16'h0739] = 8'hd0; ram[16'h073a] = 8'hfe; ram[16'h073b] = 8'h68; ram[16'h073c] = 8'h48; ram[16'h073d] = 8'hc9; ram[16'h073e] = 8'h30; ram[16'h073f] = 8'hd0; 

ram[16'h0740] = 8'hfe; ram[16'h0741] = 8'h28; ram[16'h0742] = 8'ha9; ram[16'h0743] = 8'hff; ram[16'h0744] = 8'h48; ram[16'h0745] = 8'ha9; ram[16'h0746] = 8'hcc; ram[16'h0747] = 8'h28; 
ram[16'h0748] = 8'h0f; ram[16'h0749] = 8'h0c; ram[16'h074a] = 8'h06; ram[16'h074b] = 8'h8f; ram[16'h074c] = 8'h0c; ram[16'h074d] = 8'h06; ram[16'h074e] = 8'h4c; ram[16'h074f] = 8'h4e; 
ram[16'h0750] = 8'h07; ram[16'h0751] = 8'h4c; ram[16'h0752] = 8'h51; ram[16'h0753] = 8'h07; ram[16'h0754] = 8'h08; ram[16'h0755] = 8'hc9; ram[16'h0756] = 8'hcc; ram[16'h0757] = 8'hd0; 
ram[16'h0758] = 8'hfe; ram[16'h0759] = 8'h68; ram[16'h075a] = 8'h48; ram[16'h075b] = 8'hc9; ram[16'h075c] = 8'hff; ram[16'h075d] = 8'hd0; ram[16'h075e] = 8'hfe; ram[16'h075f] = 8'h28; 

ram[16'h0760] = 8'ha5; ram[16'h0761] = 8'h0c; ram[16'h0762] = 8'hc9; ram[16'h0763] = 8'h01; ram[16'h0764] = 8'hd0; ram[16'h0765] = 8'hfe; ram[16'h0766] = 8'ha9; ram[16'h0767] = 8'hfe; 
ram[16'h0768] = 8'h85; ram[16'h0769] = 8'h0c; ram[16'h076a] = 8'ha9; ram[16'h076b] = 8'h00; ram[16'h076c] = 8'h48; ram[16'h076d] = 8'ha9; ram[16'h076e] = 8'h33; ram[16'h076f] = 8'h28; 
ram[16'h0770] = 8'h8f; ram[16'h0771] = 8'h0c; ram[16'h0772] = 8'h06; ram[16'h0773] = 8'h0f; ram[16'h0774] = 8'h0c; ram[16'h0775] = 8'h06; ram[16'h0776] = 8'h4c; ram[16'h0777] = 8'h76; 
ram[16'h0778] = 8'h07; ram[16'h0779] = 8'h4c; ram[16'h077a] = 8'h79; ram[16'h077b] = 8'h07; ram[16'h077c] = 8'h08; ram[16'h077d] = 8'hc9; ram[16'h077e] = 8'h33; ram[16'h077f] = 8'hd0; 

ram[16'h0780] = 8'hfe; ram[16'h0781] = 8'h68; ram[16'h0782] = 8'h48; ram[16'h0783] = 8'hc9; ram[16'h0784] = 8'h30; ram[16'h0785] = 8'hd0; ram[16'h0786] = 8'hfe; ram[16'h0787] = 8'h28; 
ram[16'h0788] = 8'ha9; ram[16'h0789] = 8'hff; ram[16'h078a] = 8'h48; ram[16'h078b] = 8'ha9; ram[16'h078c] = 8'hcc; ram[16'h078d] = 8'h28; ram[16'h078e] = 8'h8f; ram[16'h078f] = 8'h0c; 
ram[16'h0790] = 8'h06; ram[16'h0791] = 8'h0f; ram[16'h0792] = 8'h0c; ram[16'h0793] = 8'h06; ram[16'h0794] = 8'h4c; ram[16'h0795] = 8'h94; ram[16'h0796] = 8'h07; ram[16'h0797] = 8'h4c; 
ram[16'h0798] = 8'h97; ram[16'h0799] = 8'h07; ram[16'h079a] = 8'h08; ram[16'h079b] = 8'hc9; ram[16'h079c] = 8'hcc; ram[16'h079d] = 8'hd0; ram[16'h079e] = 8'hfe; ram[16'h079f] = 8'h68; 

ram[16'h07a0] = 8'h48; ram[16'h07a1] = 8'hc9; ram[16'h07a2] = 8'hff; ram[16'h07a3] = 8'hd0; ram[16'h07a4] = 8'hfe; ram[16'h07a5] = 8'h28; ram[16'h07a6] = 8'ha5; ram[16'h07a7] = 8'h0c; 
ram[16'h07a8] = 8'hc9; ram[16'h07a9] = 8'hfe; ram[16'h07aa] = 8'hd0; ram[16'h07ab] = 8'hfe; ram[16'h07ac] = 8'ha9; ram[16'h07ad] = 8'h02; ram[16'h07ae] = 8'h85; ram[16'h07af] = 8'h0c; 
ram[16'h07b0] = 8'ha9; ram[16'h07b1] = 8'h00; ram[16'h07b2] = 8'h48; ram[16'h07b3] = 8'ha9; ram[16'h07b4] = 8'h33; ram[16'h07b5] = 8'h28; ram[16'h07b6] = 8'h1f; ram[16'h07b7] = 8'h0c; 
ram[16'h07b8] = 8'h06; ram[16'h07b9] = 8'h9f; ram[16'h07ba] = 8'h0c; ram[16'h07bb] = 8'h06; ram[16'h07bc] = 8'h4c; ram[16'h07bd] = 8'hbc; ram[16'h07be] = 8'h07; ram[16'h07bf] = 8'h4c; 

ram[16'h07c0] = 8'hbf; ram[16'h07c1] = 8'h07; ram[16'h07c2] = 8'h08; ram[16'h07c3] = 8'hc9; ram[16'h07c4] = 8'h33; ram[16'h07c5] = 8'hd0; ram[16'h07c6] = 8'hfe; ram[16'h07c7] = 8'h68; 
ram[16'h07c8] = 8'h48; ram[16'h07c9] = 8'hc9; ram[16'h07ca] = 8'h30; ram[16'h07cb] = 8'hd0; ram[16'h07cc] = 8'hfe; ram[16'h07cd] = 8'h28; ram[16'h07ce] = 8'ha9; ram[16'h07cf] = 8'hff; 
ram[16'h07d0] = 8'h48; ram[16'h07d1] = 8'ha9; ram[16'h07d2] = 8'hcc; ram[16'h07d3] = 8'h28; ram[16'h07d4] = 8'h1f; ram[16'h07d5] = 8'h0c; ram[16'h07d6] = 8'h06; ram[16'h07d7] = 8'h9f; 
ram[16'h07d8] = 8'h0c; ram[16'h07d9] = 8'h06; ram[16'h07da] = 8'h4c; ram[16'h07db] = 8'hda; ram[16'h07dc] = 8'h07; ram[16'h07dd] = 8'h4c; ram[16'h07de] = 8'hdd; ram[16'h07df] = 8'h07; 

ram[16'h07e0] = 8'h08; ram[16'h07e1] = 8'hc9; ram[16'h07e2] = 8'hcc; ram[16'h07e3] = 8'hd0; ram[16'h07e4] = 8'hfe; ram[16'h07e5] = 8'h68; ram[16'h07e6] = 8'h48; ram[16'h07e7] = 8'hc9; 
ram[16'h07e8] = 8'hff; ram[16'h07e9] = 8'hd0; ram[16'h07ea] = 8'hfe; ram[16'h07eb] = 8'h28; ram[16'h07ec] = 8'ha5; ram[16'h07ed] = 8'h0c; ram[16'h07ee] = 8'hc9; ram[16'h07ef] = 8'h02; 
ram[16'h07f0] = 8'hd0; ram[16'h07f1] = 8'hfe; ram[16'h07f2] = 8'ha9; ram[16'h07f3] = 8'hfd; ram[16'h07f4] = 8'h85; ram[16'h07f5] = 8'h0c; ram[16'h07f6] = 8'ha9; ram[16'h07f7] = 8'h00; 
ram[16'h07f8] = 8'h48; ram[16'h07f9] = 8'ha9; ram[16'h07fa] = 8'h33; ram[16'h07fb] = 8'h28; ram[16'h07fc] = 8'h9f; ram[16'h07fd] = 8'h0c; ram[16'h07fe] = 8'h06; ram[16'h07ff] = 8'h1f; 

ram[16'h0800] = 8'h0c; ram[16'h0801] = 8'h06; ram[16'h0802] = 8'h4c; ram[16'h0803] = 8'h02; ram[16'h0804] = 8'h08; ram[16'h0805] = 8'h4c; ram[16'h0806] = 8'h05; ram[16'h0807] = 8'h08; 
ram[16'h0808] = 8'h08; ram[16'h0809] = 8'hc9; ram[16'h080a] = 8'h33; ram[16'h080b] = 8'hd0; ram[16'h080c] = 8'hfe; ram[16'h080d] = 8'h68; ram[16'h080e] = 8'h48; ram[16'h080f] = 8'hc9; 
ram[16'h0810] = 8'h30; ram[16'h0811] = 8'hd0; ram[16'h0812] = 8'hfe; ram[16'h0813] = 8'h28; ram[16'h0814] = 8'ha9; ram[16'h0815] = 8'hff; ram[16'h0816] = 8'h48; ram[16'h0817] = 8'ha9; 
ram[16'h0818] = 8'hcc; ram[16'h0819] = 8'h28; ram[16'h081a] = 8'h9f; ram[16'h081b] = 8'h0c; ram[16'h081c] = 8'h06; ram[16'h081d] = 8'h1f; ram[16'h081e] = 8'h0c; ram[16'h081f] = 8'h06; 

ram[16'h0820] = 8'h4c; ram[16'h0821] = 8'h20; ram[16'h0822] = 8'h08; ram[16'h0823] = 8'h4c; ram[16'h0824] = 8'h23; ram[16'h0825] = 8'h08; ram[16'h0826] = 8'h08; ram[16'h0827] = 8'hc9; 
ram[16'h0828] = 8'hcc; ram[16'h0829] = 8'hd0; ram[16'h082a] = 8'hfe; ram[16'h082b] = 8'h68; ram[16'h082c] = 8'h48; ram[16'h082d] = 8'hc9; ram[16'h082e] = 8'hff; ram[16'h082f] = 8'hd0; 
ram[16'h0830] = 8'hfe; ram[16'h0831] = 8'h28; ram[16'h0832] = 8'ha5; ram[16'h0833] = 8'h0c; ram[16'h0834] = 8'hc9; ram[16'h0835] = 8'hfd; ram[16'h0836] = 8'hd0; ram[16'h0837] = 8'hfe; 
ram[16'h0838] = 8'ha9; ram[16'h0839] = 8'h04; ram[16'h083a] = 8'h85; ram[16'h083b] = 8'h0c; ram[16'h083c] = 8'ha9; ram[16'h083d] = 8'h00; ram[16'h083e] = 8'h48; ram[16'h083f] = 8'ha9; 

ram[16'h0840] = 8'h33; ram[16'h0841] = 8'h28; ram[16'h0842] = 8'h2f; ram[16'h0843] = 8'h0c; ram[16'h0844] = 8'h06; ram[16'h0845] = 8'haf; ram[16'h0846] = 8'h0c; ram[16'h0847] = 8'h06; 
ram[16'h0848] = 8'h4c; ram[16'h0849] = 8'h48; ram[16'h084a] = 8'h08; ram[16'h084b] = 8'h4c; ram[16'h084c] = 8'h4b; ram[16'h084d] = 8'h08; ram[16'h084e] = 8'h08; ram[16'h084f] = 8'hc9; 
ram[16'h0850] = 8'h33; ram[16'h0851] = 8'hd0; ram[16'h0852] = 8'hfe; ram[16'h0853] = 8'h68; ram[16'h0854] = 8'h48; ram[16'h0855] = 8'hc9; ram[16'h0856] = 8'h30; ram[16'h0857] = 8'hd0; 
ram[16'h0858] = 8'hfe; ram[16'h0859] = 8'h28; ram[16'h085a] = 8'ha9; ram[16'h085b] = 8'hff; ram[16'h085c] = 8'h48; ram[16'h085d] = 8'ha9; ram[16'h085e] = 8'hcc; ram[16'h085f] = 8'h28; 

ram[16'h0860] = 8'h2f; ram[16'h0861] = 8'h0c; ram[16'h0862] = 8'h06; ram[16'h0863] = 8'haf; ram[16'h0864] = 8'h0c; ram[16'h0865] = 8'h06; ram[16'h0866] = 8'h4c; ram[16'h0867] = 8'h66; 
ram[16'h0868] = 8'h08; ram[16'h0869] = 8'h4c; ram[16'h086a] = 8'h69; ram[16'h086b] = 8'h08; ram[16'h086c] = 8'h08; ram[16'h086d] = 8'hc9; ram[16'h086e] = 8'hcc; ram[16'h086f] = 8'hd0; 
ram[16'h0870] = 8'hfe; ram[16'h0871] = 8'h68; ram[16'h0872] = 8'h48; ram[16'h0873] = 8'hc9; ram[16'h0874] = 8'hff; ram[16'h0875] = 8'hd0; ram[16'h0876] = 8'hfe; ram[16'h0877] = 8'h28; 
ram[16'h0878] = 8'ha5; ram[16'h0879] = 8'h0c; ram[16'h087a] = 8'hc9; ram[16'h087b] = 8'h04; ram[16'h087c] = 8'hd0; ram[16'h087d] = 8'hfe; ram[16'h087e] = 8'ha9; ram[16'h087f] = 8'hfb; 

ram[16'h0880] = 8'h85; ram[16'h0881] = 8'h0c; ram[16'h0882] = 8'ha9; ram[16'h0883] = 8'h00; ram[16'h0884] = 8'h48; ram[16'h0885] = 8'ha9; ram[16'h0886] = 8'h33; ram[16'h0887] = 8'h28; 
ram[16'h0888] = 8'haf; ram[16'h0889] = 8'h0c; ram[16'h088a] = 8'h06; ram[16'h088b] = 8'h2f; ram[16'h088c] = 8'h0c; ram[16'h088d] = 8'h06; ram[16'h088e] = 8'h4c; ram[16'h088f] = 8'h8e; 
ram[16'h0890] = 8'h08; ram[16'h0891] = 8'h4c; ram[16'h0892] = 8'h91; ram[16'h0893] = 8'h08; ram[16'h0894] = 8'h08; ram[16'h0895] = 8'hc9; ram[16'h0896] = 8'h33; ram[16'h0897] = 8'hd0; 
ram[16'h0898] = 8'hfe; ram[16'h0899] = 8'h68; ram[16'h089a] = 8'h48; ram[16'h089b] = 8'hc9; ram[16'h089c] = 8'h30; ram[16'h089d] = 8'hd0; ram[16'h089e] = 8'hfe; ram[16'h089f] = 8'h28; 

ram[16'h08a0] = 8'ha9; ram[16'h08a1] = 8'hff; ram[16'h08a2] = 8'h48; ram[16'h08a3] = 8'ha9; ram[16'h08a4] = 8'hcc; ram[16'h08a5] = 8'h28; ram[16'h08a6] = 8'haf; ram[16'h08a7] = 8'h0c; 
ram[16'h08a8] = 8'h06; ram[16'h08a9] = 8'h2f; ram[16'h08aa] = 8'h0c; ram[16'h08ab] = 8'h06; ram[16'h08ac] = 8'h4c; ram[16'h08ad] = 8'hac; ram[16'h08ae] = 8'h08; ram[16'h08af] = 8'h4c; 
ram[16'h08b0] = 8'haf; ram[16'h08b1] = 8'h08; ram[16'h08b2] = 8'h08; ram[16'h08b3] = 8'hc9; ram[16'h08b4] = 8'hcc; ram[16'h08b5] = 8'hd0; ram[16'h08b6] = 8'hfe; ram[16'h08b7] = 8'h68; 
ram[16'h08b8] = 8'h48; ram[16'h08b9] = 8'hc9; ram[16'h08ba] = 8'hff; ram[16'h08bb] = 8'hd0; ram[16'h08bc] = 8'hfe; ram[16'h08bd] = 8'h28; ram[16'h08be] = 8'ha5; ram[16'h08bf] = 8'h0c; 

ram[16'h08c0] = 8'hc9; ram[16'h08c1] = 8'hfb; ram[16'h08c2] = 8'hd0; ram[16'h08c3] = 8'hfe; ram[16'h08c4] = 8'ha9; ram[16'h08c5] = 8'h08; ram[16'h08c6] = 8'h85; ram[16'h08c7] = 8'h0c; 
ram[16'h08c8] = 8'ha9; ram[16'h08c9] = 8'h00; ram[16'h08ca] = 8'h48; ram[16'h08cb] = 8'ha9; ram[16'h08cc] = 8'h33; ram[16'h08cd] = 8'h28; ram[16'h08ce] = 8'h3f; ram[16'h08cf] = 8'h0c; 
ram[16'h08d0] = 8'h06; ram[16'h08d1] = 8'hbf; ram[16'h08d2] = 8'h0c; ram[16'h08d3] = 8'h06; ram[16'h08d4] = 8'h4c; ram[16'h08d5] = 8'hd4; ram[16'h08d6] = 8'h08; ram[16'h08d7] = 8'h4c; 
ram[16'h08d8] = 8'hd7; ram[16'h08d9] = 8'h08; ram[16'h08da] = 8'h08; ram[16'h08db] = 8'hc9; ram[16'h08dc] = 8'h33; ram[16'h08dd] = 8'hd0; ram[16'h08de] = 8'hfe; ram[16'h08df] = 8'h68; 

ram[16'h08e0] = 8'h48; ram[16'h08e1] = 8'hc9; ram[16'h08e2] = 8'h30; ram[16'h08e3] = 8'hd0; ram[16'h08e4] = 8'hfe; ram[16'h08e5] = 8'h28; ram[16'h08e6] = 8'ha9; ram[16'h08e7] = 8'hff; 
ram[16'h08e8] = 8'h48; ram[16'h08e9] = 8'ha9; ram[16'h08ea] = 8'hcc; ram[16'h08eb] = 8'h28; ram[16'h08ec] = 8'h3f; ram[16'h08ed] = 8'h0c; ram[16'h08ee] = 8'h06; ram[16'h08ef] = 8'hbf; 
ram[16'h08f0] = 8'h0c; ram[16'h08f1] = 8'h06; ram[16'h08f2] = 8'h4c; ram[16'h08f3] = 8'hf2; ram[16'h08f4] = 8'h08; ram[16'h08f5] = 8'h4c; ram[16'h08f6] = 8'hf5; ram[16'h08f7] = 8'h08; 
ram[16'h08f8] = 8'h08; ram[16'h08f9] = 8'hc9; ram[16'h08fa] = 8'hcc; ram[16'h08fb] = 8'hd0; ram[16'h08fc] = 8'hfe; ram[16'h08fd] = 8'h68; ram[16'h08fe] = 8'h48; ram[16'h08ff] = 8'hc9; 

ram[16'h0900] = 8'hff; ram[16'h0901] = 8'hd0; ram[16'h0902] = 8'hfe; ram[16'h0903] = 8'h28; ram[16'h0904] = 8'ha5; ram[16'h0905] = 8'h0c; ram[16'h0906] = 8'hc9; ram[16'h0907] = 8'h08; 
ram[16'h0908] = 8'hd0; ram[16'h0909] = 8'hfe; ram[16'h090a] = 8'ha9; ram[16'h090b] = 8'hf7; ram[16'h090c] = 8'h85; ram[16'h090d] = 8'h0c; ram[16'h090e] = 8'ha9; ram[16'h090f] = 8'h00; 
ram[16'h0910] = 8'h48; ram[16'h0911] = 8'ha9; ram[16'h0912] = 8'h33; ram[16'h0913] = 8'h28; ram[16'h0914] = 8'hbf; ram[16'h0915] = 8'h0c; ram[16'h0916] = 8'h06; ram[16'h0917] = 8'h3f; 
ram[16'h0918] = 8'h0c; ram[16'h0919] = 8'h06; ram[16'h091a] = 8'h4c; ram[16'h091b] = 8'h1a; ram[16'h091c] = 8'h09; ram[16'h091d] = 8'h4c; ram[16'h091e] = 8'h1d; ram[16'h091f] = 8'h09; 

ram[16'h0920] = 8'h08; ram[16'h0921] = 8'hc9; ram[16'h0922] = 8'h33; ram[16'h0923] = 8'hd0; ram[16'h0924] = 8'hfe; ram[16'h0925] = 8'h68; ram[16'h0926] = 8'h48; ram[16'h0927] = 8'hc9; 
ram[16'h0928] = 8'h30; ram[16'h0929] = 8'hd0; ram[16'h092a] = 8'hfe; ram[16'h092b] = 8'h28; ram[16'h092c] = 8'ha9; ram[16'h092d] = 8'hff; ram[16'h092e] = 8'h48; ram[16'h092f] = 8'ha9; 
ram[16'h0930] = 8'hcc; ram[16'h0931] = 8'h28; ram[16'h0932] = 8'hbf; ram[16'h0933] = 8'h0c; ram[16'h0934] = 8'h06; ram[16'h0935] = 8'h3f; ram[16'h0936] = 8'h0c; ram[16'h0937] = 8'h06; 
ram[16'h0938] = 8'h4c; ram[16'h0939] = 8'h38; ram[16'h093a] = 8'h09; ram[16'h093b] = 8'h4c; ram[16'h093c] = 8'h3b; ram[16'h093d] = 8'h09; ram[16'h093e] = 8'h08; ram[16'h093f] = 8'hc9; 

ram[16'h0940] = 8'hcc; ram[16'h0941] = 8'hd0; ram[16'h0942] = 8'hfe; ram[16'h0943] = 8'h68; ram[16'h0944] = 8'h48; ram[16'h0945] = 8'hc9; ram[16'h0946] = 8'hff; ram[16'h0947] = 8'hd0; 
ram[16'h0948] = 8'hfe; ram[16'h0949] = 8'h28; ram[16'h094a] = 8'ha5; ram[16'h094b] = 8'h0c; ram[16'h094c] = 8'hc9; ram[16'h094d] = 8'hf7; ram[16'h094e] = 8'hd0; ram[16'h094f] = 8'hfe; 
ram[16'h0950] = 8'ha9; ram[16'h0951] = 8'h10; ram[16'h0952] = 8'h85; ram[16'h0953] = 8'h0c; ram[16'h0954] = 8'ha9; ram[16'h0955] = 8'h00; ram[16'h0956] = 8'h48; ram[16'h0957] = 8'ha9; 
ram[16'h0958] = 8'h33; ram[16'h0959] = 8'h28; ram[16'h095a] = 8'h4f; ram[16'h095b] = 8'h0c; ram[16'h095c] = 8'h06; ram[16'h095d] = 8'hcf; ram[16'h095e] = 8'h0c; ram[16'h095f] = 8'h06; 

ram[16'h0960] = 8'h4c; ram[16'h0961] = 8'h60; ram[16'h0962] = 8'h09; ram[16'h0963] = 8'h4c; ram[16'h0964] = 8'h63; ram[16'h0965] = 8'h09; ram[16'h0966] = 8'h08; ram[16'h0967] = 8'hc9; 
ram[16'h0968] = 8'h33; ram[16'h0969] = 8'hd0; ram[16'h096a] = 8'hfe; ram[16'h096b] = 8'h68; ram[16'h096c] = 8'h48; ram[16'h096d] = 8'hc9; ram[16'h096e] = 8'h30; ram[16'h096f] = 8'hd0; 
ram[16'h0970] = 8'hfe; ram[16'h0971] = 8'h28; ram[16'h0972] = 8'ha9; ram[16'h0973] = 8'hff; ram[16'h0974] = 8'h48; ram[16'h0975] = 8'ha9; ram[16'h0976] = 8'hcc; ram[16'h0977] = 8'h28; 
ram[16'h0978] = 8'h4f; ram[16'h0979] = 8'h0c; ram[16'h097a] = 8'h06; ram[16'h097b] = 8'hcf; ram[16'h097c] = 8'h0c; ram[16'h097d] = 8'h06; ram[16'h097e] = 8'h4c; ram[16'h097f] = 8'h7e; 

ram[16'h0980] = 8'h09; ram[16'h0981] = 8'h4c; ram[16'h0982] = 8'h81; ram[16'h0983] = 8'h09; ram[16'h0984] = 8'h08; ram[16'h0985] = 8'hc9; ram[16'h0986] = 8'hcc; ram[16'h0987] = 8'hd0; 
ram[16'h0988] = 8'hfe; ram[16'h0989] = 8'h68; ram[16'h098a] = 8'h48; ram[16'h098b] = 8'hc9; ram[16'h098c] = 8'hff; ram[16'h098d] = 8'hd0; ram[16'h098e] = 8'hfe; ram[16'h098f] = 8'h28; 
ram[16'h0990] = 8'ha5; ram[16'h0991] = 8'h0c; ram[16'h0992] = 8'hc9; ram[16'h0993] = 8'h10; ram[16'h0994] = 8'hd0; ram[16'h0995] = 8'hfe; ram[16'h0996] = 8'ha9; ram[16'h0997] = 8'hef; 
ram[16'h0998] = 8'h85; ram[16'h0999] = 8'h0c; ram[16'h099a] = 8'ha9; ram[16'h099b] = 8'h00; ram[16'h099c] = 8'h48; ram[16'h099d] = 8'ha9; ram[16'h099e] = 8'h33; ram[16'h099f] = 8'h28; 

ram[16'h09a0] = 8'hcf; ram[16'h09a1] = 8'h0c; ram[16'h09a2] = 8'h06; ram[16'h09a3] = 8'h4f; ram[16'h09a4] = 8'h0c; ram[16'h09a5] = 8'h06; ram[16'h09a6] = 8'h4c; ram[16'h09a7] = 8'ha6; 
ram[16'h09a8] = 8'h09; ram[16'h09a9] = 8'h4c; ram[16'h09aa] = 8'ha9; ram[16'h09ab] = 8'h09; ram[16'h09ac] = 8'h08; ram[16'h09ad] = 8'hc9; ram[16'h09ae] = 8'h33; ram[16'h09af] = 8'hd0; 
ram[16'h09b0] = 8'hfe; ram[16'h09b1] = 8'h68; ram[16'h09b2] = 8'h48; ram[16'h09b3] = 8'hc9; ram[16'h09b4] = 8'h30; ram[16'h09b5] = 8'hd0; ram[16'h09b6] = 8'hfe; ram[16'h09b7] = 8'h28; 
ram[16'h09b8] = 8'ha9; ram[16'h09b9] = 8'hff; ram[16'h09ba] = 8'h48; ram[16'h09bb] = 8'ha9; ram[16'h09bc] = 8'hcc; ram[16'h09bd] = 8'h28; ram[16'h09be] = 8'hcf; ram[16'h09bf] = 8'h0c; 

ram[16'h09c0] = 8'h06; ram[16'h09c1] = 8'h4f; ram[16'h09c2] = 8'h0c; ram[16'h09c3] = 8'h06; ram[16'h09c4] = 8'h4c; ram[16'h09c5] = 8'hc4; ram[16'h09c6] = 8'h09; ram[16'h09c7] = 8'h4c; 
ram[16'h09c8] = 8'hc7; ram[16'h09c9] = 8'h09; ram[16'h09ca] = 8'h08; ram[16'h09cb] = 8'hc9; ram[16'h09cc] = 8'hcc; ram[16'h09cd] = 8'hd0; ram[16'h09ce] = 8'hfe; ram[16'h09cf] = 8'h68; 
ram[16'h09d0] = 8'h48; ram[16'h09d1] = 8'hc9; ram[16'h09d2] = 8'hff; ram[16'h09d3] = 8'hd0; ram[16'h09d4] = 8'hfe; ram[16'h09d5] = 8'h28; ram[16'h09d6] = 8'ha5; ram[16'h09d7] = 8'h0c; 
ram[16'h09d8] = 8'hc9; ram[16'h09d9] = 8'hef; ram[16'h09da] = 8'hd0; ram[16'h09db] = 8'hfe; ram[16'h09dc] = 8'ha9; ram[16'h09dd] = 8'h20; ram[16'h09de] = 8'h85; ram[16'h09df] = 8'h0c; 

ram[16'h09e0] = 8'ha9; ram[16'h09e1] = 8'h00; ram[16'h09e2] = 8'h48; ram[16'h09e3] = 8'ha9; ram[16'h09e4] = 8'h33; ram[16'h09e5] = 8'h28; ram[16'h09e6] = 8'h5f; ram[16'h09e7] = 8'h0c; 
ram[16'h09e8] = 8'h06; ram[16'h09e9] = 8'hdf; ram[16'h09ea] = 8'h0c; ram[16'h09eb] = 8'h06; ram[16'h09ec] = 8'h4c; ram[16'h09ed] = 8'hec; ram[16'h09ee] = 8'h09; ram[16'h09ef] = 8'h4c; 
ram[16'h09f0] = 8'hef; ram[16'h09f1] = 8'h09; ram[16'h09f2] = 8'h08; ram[16'h09f3] = 8'hc9; ram[16'h09f4] = 8'h33; ram[16'h09f5] = 8'hd0; ram[16'h09f6] = 8'hfe; ram[16'h09f7] = 8'h68; 
ram[16'h09f8] = 8'h48; ram[16'h09f9] = 8'hc9; ram[16'h09fa] = 8'h30; ram[16'h09fb] = 8'hd0; ram[16'h09fc] = 8'hfe; ram[16'h09fd] = 8'h28; ram[16'h09fe] = 8'ha9; ram[16'h09ff] = 8'hff; 

ram[16'h0a00] = 8'h48; ram[16'h0a01] = 8'ha9; ram[16'h0a02] = 8'hcc; ram[16'h0a03] = 8'h28; ram[16'h0a04] = 8'h5f; ram[16'h0a05] = 8'h0c; ram[16'h0a06] = 8'h06; ram[16'h0a07] = 8'hdf; 
ram[16'h0a08] = 8'h0c; ram[16'h0a09] = 8'h06; ram[16'h0a0a] = 8'h4c; ram[16'h0a0b] = 8'h0a; ram[16'h0a0c] = 8'h0a; ram[16'h0a0d] = 8'h4c; ram[16'h0a0e] = 8'h0d; ram[16'h0a0f] = 8'h0a; 
ram[16'h0a10] = 8'h08; ram[16'h0a11] = 8'hc9; ram[16'h0a12] = 8'hcc; ram[16'h0a13] = 8'hd0; ram[16'h0a14] = 8'hfe; ram[16'h0a15] = 8'h68; ram[16'h0a16] = 8'h48; ram[16'h0a17] = 8'hc9; 
ram[16'h0a18] = 8'hff; ram[16'h0a19] = 8'hd0; ram[16'h0a1a] = 8'hfe; ram[16'h0a1b] = 8'h28; ram[16'h0a1c] = 8'ha5; ram[16'h0a1d] = 8'h0c; ram[16'h0a1e] = 8'hc9; ram[16'h0a1f] = 8'h20; 

ram[16'h0a20] = 8'hd0; ram[16'h0a21] = 8'hfe; ram[16'h0a22] = 8'ha9; ram[16'h0a23] = 8'hdf; ram[16'h0a24] = 8'h85; ram[16'h0a25] = 8'h0c; ram[16'h0a26] = 8'ha9; ram[16'h0a27] = 8'h00; 
ram[16'h0a28] = 8'h48; ram[16'h0a29] = 8'ha9; ram[16'h0a2a] = 8'h33; ram[16'h0a2b] = 8'h28; ram[16'h0a2c] = 8'hdf; ram[16'h0a2d] = 8'h0c; ram[16'h0a2e] = 8'h06; ram[16'h0a2f] = 8'h5f; 
ram[16'h0a30] = 8'h0c; ram[16'h0a31] = 8'h06; ram[16'h0a32] = 8'h4c; ram[16'h0a33] = 8'h32; ram[16'h0a34] = 8'h0a; ram[16'h0a35] = 8'h4c; ram[16'h0a36] = 8'h35; ram[16'h0a37] = 8'h0a; 
ram[16'h0a38] = 8'h08; ram[16'h0a39] = 8'hc9; ram[16'h0a3a] = 8'h33; ram[16'h0a3b] = 8'hd0; ram[16'h0a3c] = 8'hfe; ram[16'h0a3d] = 8'h68; ram[16'h0a3e] = 8'h48; ram[16'h0a3f] = 8'hc9; 

ram[16'h0a40] = 8'h30; ram[16'h0a41] = 8'hd0; ram[16'h0a42] = 8'hfe; ram[16'h0a43] = 8'h28; ram[16'h0a44] = 8'ha9; ram[16'h0a45] = 8'hff; ram[16'h0a46] = 8'h48; ram[16'h0a47] = 8'ha9; 
ram[16'h0a48] = 8'hcc; ram[16'h0a49] = 8'h28; ram[16'h0a4a] = 8'hdf; ram[16'h0a4b] = 8'h0c; ram[16'h0a4c] = 8'h06; ram[16'h0a4d] = 8'h5f; ram[16'h0a4e] = 8'h0c; ram[16'h0a4f] = 8'h06; 
ram[16'h0a50] = 8'h4c; ram[16'h0a51] = 8'h50; ram[16'h0a52] = 8'h0a; ram[16'h0a53] = 8'h4c; ram[16'h0a54] = 8'h53; ram[16'h0a55] = 8'h0a; ram[16'h0a56] = 8'h08; ram[16'h0a57] = 8'hc9; 
ram[16'h0a58] = 8'hcc; ram[16'h0a59] = 8'hd0; ram[16'h0a5a] = 8'hfe; ram[16'h0a5b] = 8'h68; ram[16'h0a5c] = 8'h48; ram[16'h0a5d] = 8'hc9; ram[16'h0a5e] = 8'hff; ram[16'h0a5f] = 8'hd0; 

ram[16'h0a60] = 8'hfe; ram[16'h0a61] = 8'h28; ram[16'h0a62] = 8'ha5; ram[16'h0a63] = 8'h0c; ram[16'h0a64] = 8'hc9; ram[16'h0a65] = 8'hdf; ram[16'h0a66] = 8'hd0; ram[16'h0a67] = 8'hfe; 
ram[16'h0a68] = 8'ha9; ram[16'h0a69] = 8'h40; ram[16'h0a6a] = 8'h85; ram[16'h0a6b] = 8'h0c; ram[16'h0a6c] = 8'ha9; ram[16'h0a6d] = 8'h00; ram[16'h0a6e] = 8'h48; ram[16'h0a6f] = 8'ha9; 
ram[16'h0a70] = 8'h33; ram[16'h0a71] = 8'h28; ram[16'h0a72] = 8'h6f; ram[16'h0a73] = 8'h0c; ram[16'h0a74] = 8'h06; ram[16'h0a75] = 8'hef; ram[16'h0a76] = 8'h0c; ram[16'h0a77] = 8'h06; 
ram[16'h0a78] = 8'h4c; ram[16'h0a79] = 8'h78; ram[16'h0a7a] = 8'h0a; ram[16'h0a7b] = 8'h4c; ram[16'h0a7c] = 8'h7b; ram[16'h0a7d] = 8'h0a; ram[16'h0a7e] = 8'h08; ram[16'h0a7f] = 8'hc9; 

ram[16'h0a80] = 8'h33; ram[16'h0a81] = 8'hd0; ram[16'h0a82] = 8'hfe; ram[16'h0a83] = 8'h68; ram[16'h0a84] = 8'h48; ram[16'h0a85] = 8'hc9; ram[16'h0a86] = 8'h30; ram[16'h0a87] = 8'hd0; 
ram[16'h0a88] = 8'hfe; ram[16'h0a89] = 8'h28; ram[16'h0a8a] = 8'ha9; ram[16'h0a8b] = 8'hff; ram[16'h0a8c] = 8'h48; ram[16'h0a8d] = 8'ha9; ram[16'h0a8e] = 8'hcc; ram[16'h0a8f] = 8'h28; 
ram[16'h0a90] = 8'h6f; ram[16'h0a91] = 8'h0c; ram[16'h0a92] = 8'h06; ram[16'h0a93] = 8'hef; ram[16'h0a94] = 8'h0c; ram[16'h0a95] = 8'h06; ram[16'h0a96] = 8'h4c; ram[16'h0a97] = 8'h96; 
ram[16'h0a98] = 8'h0a; ram[16'h0a99] = 8'h4c; ram[16'h0a9a] = 8'h99; ram[16'h0a9b] = 8'h0a; ram[16'h0a9c] = 8'h08; ram[16'h0a9d] = 8'hc9; ram[16'h0a9e] = 8'hcc; ram[16'h0a9f] = 8'hd0; 

ram[16'h0aa0] = 8'hfe; ram[16'h0aa1] = 8'h68; ram[16'h0aa2] = 8'h48; ram[16'h0aa3] = 8'hc9; ram[16'h0aa4] = 8'hff; ram[16'h0aa5] = 8'hd0; ram[16'h0aa6] = 8'hfe; ram[16'h0aa7] = 8'h28; 
ram[16'h0aa8] = 8'ha5; ram[16'h0aa9] = 8'h0c; ram[16'h0aaa] = 8'hc9; ram[16'h0aab] = 8'h40; ram[16'h0aac] = 8'hd0; ram[16'h0aad] = 8'hfe; ram[16'h0aae] = 8'ha9; ram[16'h0aaf] = 8'hbf; 
ram[16'h0ab0] = 8'h85; ram[16'h0ab1] = 8'h0c; ram[16'h0ab2] = 8'ha9; ram[16'h0ab3] = 8'h00; ram[16'h0ab4] = 8'h48; ram[16'h0ab5] = 8'ha9; ram[16'h0ab6] = 8'h33; ram[16'h0ab7] = 8'h28; 
ram[16'h0ab8] = 8'hef; ram[16'h0ab9] = 8'h0c; ram[16'h0aba] = 8'h06; ram[16'h0abb] = 8'h6f; ram[16'h0abc] = 8'h0c; ram[16'h0abd] = 8'h06; ram[16'h0abe] = 8'h4c; ram[16'h0abf] = 8'hbe; 

ram[16'h0ac0] = 8'h0a; ram[16'h0ac1] = 8'h4c; ram[16'h0ac2] = 8'hc1; ram[16'h0ac3] = 8'h0a; ram[16'h0ac4] = 8'h08; ram[16'h0ac5] = 8'hc9; ram[16'h0ac6] = 8'h33; ram[16'h0ac7] = 8'hd0; 
ram[16'h0ac8] = 8'hfe; ram[16'h0ac9] = 8'h68; ram[16'h0aca] = 8'h48; ram[16'h0acb] = 8'hc9; ram[16'h0acc] = 8'h30; ram[16'h0acd] = 8'hd0; ram[16'h0ace] = 8'hfe; ram[16'h0acf] = 8'h28; 
ram[16'h0ad0] = 8'ha9; ram[16'h0ad1] = 8'hff; ram[16'h0ad2] = 8'h48; ram[16'h0ad3] = 8'ha9; ram[16'h0ad4] = 8'hcc; ram[16'h0ad5] = 8'h28; ram[16'h0ad6] = 8'hef; ram[16'h0ad7] = 8'h0c; 
ram[16'h0ad8] = 8'h06; ram[16'h0ad9] = 8'h6f; ram[16'h0ada] = 8'h0c; ram[16'h0adb] = 8'h06; ram[16'h0adc] = 8'h4c; ram[16'h0add] = 8'hdc; ram[16'h0ade] = 8'h0a; ram[16'h0adf] = 8'h4c; 

ram[16'h0ae0] = 8'hdf; ram[16'h0ae1] = 8'h0a; ram[16'h0ae2] = 8'h08; ram[16'h0ae3] = 8'hc9; ram[16'h0ae4] = 8'hcc; ram[16'h0ae5] = 8'hd0; ram[16'h0ae6] = 8'hfe; ram[16'h0ae7] = 8'h68; 
ram[16'h0ae8] = 8'h48; ram[16'h0ae9] = 8'hc9; ram[16'h0aea] = 8'hff; ram[16'h0aeb] = 8'hd0; ram[16'h0aec] = 8'hfe; ram[16'h0aed] = 8'h28; ram[16'h0aee] = 8'ha5; ram[16'h0aef] = 8'h0c; 
ram[16'h0af0] = 8'hc9; ram[16'h0af1] = 8'hbf; ram[16'h0af2] = 8'hd0; ram[16'h0af3] = 8'hfe; ram[16'h0af4] = 8'ha9; ram[16'h0af5] = 8'h80; ram[16'h0af6] = 8'h85; ram[16'h0af7] = 8'h0c; 
ram[16'h0af8] = 8'ha9; ram[16'h0af9] = 8'h00; ram[16'h0afa] = 8'h48; ram[16'h0afb] = 8'ha9; ram[16'h0afc] = 8'h33; ram[16'h0afd] = 8'h28; ram[16'h0afe] = 8'h7f; ram[16'h0aff] = 8'h0c; 

ram[16'h0b00] = 8'h06; ram[16'h0b01] = 8'hff; ram[16'h0b02] = 8'h0c; ram[16'h0b03] = 8'h06; ram[16'h0b04] = 8'h4c; ram[16'h0b05] = 8'h04; ram[16'h0b06] = 8'h0b; ram[16'h0b07] = 8'h4c; 
ram[16'h0b08] = 8'h07; ram[16'h0b09] = 8'h0b; ram[16'h0b0a] = 8'h08; ram[16'h0b0b] = 8'hc9; ram[16'h0b0c] = 8'h33; ram[16'h0b0d] = 8'hd0; ram[16'h0b0e] = 8'hfe; ram[16'h0b0f] = 8'h68; 
ram[16'h0b10] = 8'h48; ram[16'h0b11] = 8'hc9; ram[16'h0b12] = 8'h30; ram[16'h0b13] = 8'hd0; ram[16'h0b14] = 8'hfe; ram[16'h0b15] = 8'h28; ram[16'h0b16] = 8'ha9; ram[16'h0b17] = 8'hff; 
ram[16'h0b18] = 8'h48; ram[16'h0b19] = 8'ha9; ram[16'h0b1a] = 8'hcc; ram[16'h0b1b] = 8'h28; ram[16'h0b1c] = 8'h7f; ram[16'h0b1d] = 8'h0c; ram[16'h0b1e] = 8'h06; ram[16'h0b1f] = 8'hff; 

ram[16'h0b20] = 8'h0c; ram[16'h0b21] = 8'h06; ram[16'h0b22] = 8'h4c; ram[16'h0b23] = 8'h22; ram[16'h0b24] = 8'h0b; ram[16'h0b25] = 8'h4c; ram[16'h0b26] = 8'h25; ram[16'h0b27] = 8'h0b; 
ram[16'h0b28] = 8'h08; ram[16'h0b29] = 8'hc9; ram[16'h0b2a] = 8'hcc; ram[16'h0b2b] = 8'hd0; ram[16'h0b2c] = 8'hfe; ram[16'h0b2d] = 8'h68; ram[16'h0b2e] = 8'h48; ram[16'h0b2f] = 8'hc9; 
ram[16'h0b30] = 8'hff; ram[16'h0b31] = 8'hd0; ram[16'h0b32] = 8'hfe; ram[16'h0b33] = 8'h28; ram[16'h0b34] = 8'ha5; ram[16'h0b35] = 8'h0c; ram[16'h0b36] = 8'hc9; ram[16'h0b37] = 8'h80; 
ram[16'h0b38] = 8'hd0; ram[16'h0b39] = 8'hfe; ram[16'h0b3a] = 8'ha9; ram[16'h0b3b] = 8'h7f; ram[16'h0b3c] = 8'h85; ram[16'h0b3d] = 8'h0c; ram[16'h0b3e] = 8'ha9; ram[16'h0b3f] = 8'h00; 

ram[16'h0b40] = 8'h48; ram[16'h0b41] = 8'ha9; ram[16'h0b42] = 8'h33; ram[16'h0b43] = 8'h28; ram[16'h0b44] = 8'hff; ram[16'h0b45] = 8'h0c; ram[16'h0b46] = 8'h06; ram[16'h0b47] = 8'h7f; 
ram[16'h0b48] = 8'h0c; ram[16'h0b49] = 8'h06; ram[16'h0b4a] = 8'h4c; ram[16'h0b4b] = 8'h4a; ram[16'h0b4c] = 8'h0b; ram[16'h0b4d] = 8'h4c; ram[16'h0b4e] = 8'h4d; ram[16'h0b4f] = 8'h0b; 
ram[16'h0b50] = 8'h08; ram[16'h0b51] = 8'hc9; ram[16'h0b52] = 8'h33; ram[16'h0b53] = 8'hd0; ram[16'h0b54] = 8'hfe; ram[16'h0b55] = 8'h68; ram[16'h0b56] = 8'h48; ram[16'h0b57] = 8'hc9; 
ram[16'h0b58] = 8'h30; ram[16'h0b59] = 8'hd0; ram[16'h0b5a] = 8'hfe; ram[16'h0b5b] = 8'h28; ram[16'h0b5c] = 8'ha9; ram[16'h0b5d] = 8'hff; ram[16'h0b5e] = 8'h48; ram[16'h0b5f] = 8'ha9; 

ram[16'h0b60] = 8'hcc; ram[16'h0b61] = 8'h28; ram[16'h0b62] = 8'hff; ram[16'h0b63] = 8'h0c; ram[16'h0b64] = 8'h06; ram[16'h0b65] = 8'h7f; ram[16'h0b66] = 8'h0c; ram[16'h0b67] = 8'h06; 
ram[16'h0b68] = 8'h4c; ram[16'h0b69] = 8'h68; ram[16'h0b6a] = 8'h0b; ram[16'h0b6b] = 8'h4c; ram[16'h0b6c] = 8'h6b; ram[16'h0b6d] = 8'h0b; ram[16'h0b6e] = 8'h08; ram[16'h0b6f] = 8'hc9; 
ram[16'h0b70] = 8'hcc; ram[16'h0b71] = 8'hd0; ram[16'h0b72] = 8'hfe; ram[16'h0b73] = 8'h68; ram[16'h0b74] = 8'h48; ram[16'h0b75] = 8'hc9; ram[16'h0b76] = 8'hff; ram[16'h0b77] = 8'hd0; 
ram[16'h0b78] = 8'hfe; ram[16'h0b79] = 8'h28; ram[16'h0b7a] = 8'ha5; ram[16'h0b7b] = 8'h0c; ram[16'h0b7c] = 8'hc9; ram[16'h0b7d] = 8'h7f; ram[16'h0b7e] = 8'hd0; ram[16'h0b7f] = 8'hfe; 

ram[16'h0b80] = 8'he0; ram[16'h0b81] = 8'h11; ram[16'h0b82] = 8'hd0; ram[16'h0b83] = 8'hfe; ram[16'h0b84] = 8'hc0; ram[16'h0b85] = 8'h22; ram[16'h0b86] = 8'hd0; ram[16'h0b87] = 8'hfe; 
ram[16'h0b88] = 8'had; ram[16'h0b89] = 8'h02; ram[16'h0b8a] = 8'h02; ram[16'h0b8b] = 8'hc9; ram[16'h0b8c] = 8'h06; ram[16'h0b8d] = 8'hd0; ram[16'h0b8e] = 8'hfe; ram[16'h0b8f] = 8'ha9; 
ram[16'h0b90] = 8'h07; ram[16'h0b91] = 8'h8d; ram[16'h0b92] = 8'h02; ram[16'h0b93] = 8'h02; ram[16'h0b94] = 8'ha9; ram[16'h0b95] = 8'h00; ram[16'h0b96] = 8'h85; ram[16'h0b97] = 8'h0c; 
ram[16'h0b98] = 8'ha9; ram[16'h0b99] = 8'h00; ram[16'h0b9a] = 8'h0f; ram[16'h0b9b] = 8'h0c; ram[16'h0b9c] = 8'h02; ram[16'h0b9d] = 8'h49; ram[16'h0b9e] = 8'h01; ram[16'h0b9f] = 8'h1f; 

ram[16'h0ba0] = 8'h0c; ram[16'h0ba1] = 8'h02; ram[16'h0ba2] = 8'h49; ram[16'h0ba3] = 8'h02; ram[16'h0ba4] = 8'h2f; ram[16'h0ba5] = 8'h0c; ram[16'h0ba6] = 8'h02; ram[16'h0ba7] = 8'h49; 
ram[16'h0ba8] = 8'h04; ram[16'h0ba9] = 8'h3f; ram[16'h0baa] = 8'h0c; ram[16'h0bab] = 8'h02; ram[16'h0bac] = 8'h49; ram[16'h0bad] = 8'h08; ram[16'h0bae] = 8'h4f; ram[16'h0baf] = 8'h0c; 
ram[16'h0bb0] = 8'h02; ram[16'h0bb1] = 8'h49; ram[16'h0bb2] = 8'h10; ram[16'h0bb3] = 8'h5f; ram[16'h0bb4] = 8'h0c; ram[16'h0bb5] = 8'h02; ram[16'h0bb6] = 8'h49; ram[16'h0bb7] = 8'h20; 
ram[16'h0bb8] = 8'h6f; ram[16'h0bb9] = 8'h0c; ram[16'h0bba] = 8'h02; ram[16'h0bbb] = 8'h49; ram[16'h0bbc] = 8'h40; ram[16'h0bbd] = 8'h7f; ram[16'h0bbe] = 8'h0c; ram[16'h0bbf] = 8'h02; 

ram[16'h0bc0] = 8'h49; ram[16'h0bc1] = 8'h80; ram[16'h0bc2] = 8'h45; ram[16'h0bc3] = 8'h0c; ram[16'h0bc4] = 8'hd0; ram[16'h0bc5] = 8'hfe; ram[16'h0bc6] = 8'ha9; ram[16'h0bc7] = 8'hff; 
ram[16'h0bc8] = 8'h8f; ram[16'h0bc9] = 8'h0c; ram[16'h0bca] = 8'h02; ram[16'h0bcb] = 8'h49; ram[16'h0bcc] = 8'h01; ram[16'h0bcd] = 8'h9f; ram[16'h0bce] = 8'h0c; ram[16'h0bcf] = 8'h02; 
ram[16'h0bd0] = 8'h49; ram[16'h0bd1] = 8'h02; ram[16'h0bd2] = 8'haf; ram[16'h0bd3] = 8'h0c; ram[16'h0bd4] = 8'h02; ram[16'h0bd5] = 8'h49; ram[16'h0bd6] = 8'h04; ram[16'h0bd7] = 8'hbf; 
ram[16'h0bd8] = 8'h0c; ram[16'h0bd9] = 8'h02; ram[16'h0bda] = 8'h49; ram[16'h0bdb] = 8'h08; ram[16'h0bdc] = 8'hcf; ram[16'h0bdd] = 8'h0c; ram[16'h0bde] = 8'h02; ram[16'h0bdf] = 8'h49; 

ram[16'h0be0] = 8'h10; ram[16'h0be1] = 8'hdf; ram[16'h0be2] = 8'h0c; ram[16'h0be3] = 8'h02; ram[16'h0be4] = 8'h49; ram[16'h0be5] = 8'h20; ram[16'h0be6] = 8'hef; ram[16'h0be7] = 8'h0c; 
ram[16'h0be8] = 8'h02; ram[16'h0be9] = 8'h49; ram[16'h0bea] = 8'h40; ram[16'h0beb] = 8'hff; ram[16'h0bec] = 8'h0c; ram[16'h0bed] = 8'h02; ram[16'h0bee] = 8'h49; ram[16'h0bef] = 8'h80; 
ram[16'h0bf0] = 8'h45; ram[16'h0bf1] = 8'h0c; ram[16'h0bf2] = 8'hd0; ram[16'h0bf3] = 8'hfe; ram[16'h0bf4] = 8'he6; ram[16'h0bf5] = 8'h0c; ram[16'h0bf6] = 8'hd0; ram[16'h0bf7] = 8'ha0; 
ram[16'h0bf8] = 8'had; ram[16'h0bf9] = 8'h02; ram[16'h0bfa] = 8'h02; ram[16'h0bfb] = 8'hc9; ram[16'h0bfc] = 8'h07; ram[16'h0bfd] = 8'hd0; ram[16'h0bfe] = 8'hfe; ram[16'h0bff] = 8'ha9; 

ram[16'h0c00] = 8'h08; ram[16'h0c01] = 8'h8d; ram[16'h0c02] = 8'h02; ram[16'h0c03] = 8'h02; ram[16'h0c04] = 8'ha0; ram[16'h0c05] = 8'h42; ram[16'h0c06] = 8'ha2; ram[16'h0c07] = 8'h02; 
ram[16'h0c08] = 8'h02; ram[16'h0c09] = 8'hc8; ram[16'h0c0a] = 8'hca; ram[16'h0c0b] = 8'hca; ram[16'h0c0c] = 8'hd0; ram[16'h0c0d] = 8'hfe; ram[16'h0c0e] = 8'ha9; ram[16'h0c0f] = 8'h00; 
ram[16'h0c10] = 8'h48; ram[16'h0c11] = 8'ha9; ram[16'h0c12] = 8'hfd; ram[16'h0c13] = 8'h28; ram[16'h0c14] = 8'h02; ram[16'h0c15] = 8'hea; ram[16'h0c16] = 8'hea; ram[16'h0c17] = 8'h08; 
ram[16'h0c18] = 8'hc9; ram[16'h0c19] = 8'hfd; ram[16'h0c1a] = 8'hd0; ram[16'h0c1b] = 8'hfe; ram[16'h0c1c] = 8'h68; ram[16'h0c1d] = 8'h48; ram[16'h0c1e] = 8'hc9; ram[16'h0c1f] = 8'h30; 

ram[16'h0c20] = 8'hd0; ram[16'h0c21] = 8'hfe; ram[16'h0c22] = 8'h28; ram[16'h0c23] = 8'ha9; ram[16'h0c24] = 8'hff; ram[16'h0c25] = 8'h48; ram[16'h0c26] = 8'ha9; ram[16'h0c27] = 8'ha8; 
ram[16'h0c28] = 8'h28; ram[16'h0c29] = 8'h02; ram[16'h0c2a] = 8'hea; ram[16'h0c2b] = 8'hea; ram[16'h0c2c] = 8'h08; ram[16'h0c2d] = 8'hc9; ram[16'h0c2e] = 8'ha8; ram[16'h0c2f] = 8'hd0; 
ram[16'h0c30] = 8'hfe; ram[16'h0c31] = 8'h68; ram[16'h0c32] = 8'h48; ram[16'h0c33] = 8'hc9; ram[16'h0c34] = 8'hff; ram[16'h0c35] = 8'hd0; ram[16'h0c36] = 8'hfe; ram[16'h0c37] = 8'h28; 
ram[16'h0c38] = 8'hc0; ram[16'h0c39] = 8'h42; ram[16'h0c3a] = 8'hd0; ram[16'h0c3b] = 8'hfe; ram[16'h0c3c] = 8'he0; ram[16'h0c3d] = 8'h00; ram[16'h0c3e] = 8'hd0; ram[16'h0c3f] = 8'hfe; 

ram[16'h0c40] = 8'ha0; ram[16'h0c41] = 8'h42; ram[16'h0c42] = 8'ha2; ram[16'h0c43] = 8'h02; ram[16'h0c44] = 8'h22; ram[16'h0c45] = 8'hc8; ram[16'h0c46] = 8'hca; ram[16'h0c47] = 8'hca; 
ram[16'h0c48] = 8'hd0; ram[16'h0c49] = 8'hfe; ram[16'h0c4a] = 8'ha9; ram[16'h0c4b] = 8'h00; ram[16'h0c4c] = 8'h48; ram[16'h0c4d] = 8'ha9; ram[16'h0c4e] = 8'hdd; ram[16'h0c4f] = 8'h28; 
ram[16'h0c50] = 8'h22; ram[16'h0c51] = 8'hea; ram[16'h0c52] = 8'hea; ram[16'h0c53] = 8'h08; ram[16'h0c54] = 8'hc9; ram[16'h0c55] = 8'hdd; ram[16'h0c56] = 8'hd0; ram[16'h0c57] = 8'hfe; 
ram[16'h0c58] = 8'h68; ram[16'h0c59] = 8'h48; ram[16'h0c5a] = 8'hc9; ram[16'h0c5b] = 8'h30; ram[16'h0c5c] = 8'hd0; ram[16'h0c5d] = 8'hfe; ram[16'h0c5e] = 8'h28; ram[16'h0c5f] = 8'ha9; 

ram[16'h0c60] = 8'hff; ram[16'h0c61] = 8'h48; ram[16'h0c62] = 8'ha9; ram[16'h0c63] = 8'h88; ram[16'h0c64] = 8'h28; ram[16'h0c65] = 8'h22; ram[16'h0c66] = 8'hea; ram[16'h0c67] = 8'hea; 
ram[16'h0c68] = 8'h08; ram[16'h0c69] = 8'hc9; ram[16'h0c6a] = 8'h88; ram[16'h0c6b] = 8'hd0; ram[16'h0c6c] = 8'hfe; ram[16'h0c6d] = 8'h68; ram[16'h0c6e] = 8'h48; ram[16'h0c6f] = 8'hc9; 
ram[16'h0c70] = 8'hff; ram[16'h0c71] = 8'hd0; ram[16'h0c72] = 8'hfe; ram[16'h0c73] = 8'h28; ram[16'h0c74] = 8'hc0; ram[16'h0c75] = 8'h42; ram[16'h0c76] = 8'hd0; ram[16'h0c77] = 8'hfe; 
ram[16'h0c78] = 8'he0; ram[16'h0c79] = 8'h00; ram[16'h0c7a] = 8'hd0; ram[16'h0c7b] = 8'hfe; ram[16'h0c7c] = 8'ha0; ram[16'h0c7d] = 8'h42; ram[16'h0c7e] = 8'ha2; ram[16'h0c7f] = 8'h02; 

ram[16'h0c80] = 8'h42; ram[16'h0c81] = 8'hc8; ram[16'h0c82] = 8'hca; ram[16'h0c83] = 8'hca; ram[16'h0c84] = 8'hd0; ram[16'h0c85] = 8'hfe; ram[16'h0c86] = 8'ha9; ram[16'h0c87] = 8'h00; 
ram[16'h0c88] = 8'h48; ram[16'h0c89] = 8'ha9; ram[16'h0c8a] = 8'hbd; ram[16'h0c8b] = 8'h28; ram[16'h0c8c] = 8'h42; ram[16'h0c8d] = 8'hea; ram[16'h0c8e] = 8'hea; ram[16'h0c8f] = 8'h08; 
ram[16'h0c90] = 8'hc9; ram[16'h0c91] = 8'hbd; ram[16'h0c92] = 8'hd0; ram[16'h0c93] = 8'hfe; ram[16'h0c94] = 8'h68; ram[16'h0c95] = 8'h48; ram[16'h0c96] = 8'hc9; ram[16'h0c97] = 8'h30; 
ram[16'h0c98] = 8'hd0; ram[16'h0c99] = 8'hfe; ram[16'h0c9a] = 8'h28; ram[16'h0c9b] = 8'ha9; ram[16'h0c9c] = 8'hff; ram[16'h0c9d] = 8'h48; ram[16'h0c9e] = 8'ha9; ram[16'h0c9f] = 8'h68; 

ram[16'h0ca0] = 8'h28; ram[16'h0ca1] = 8'h42; ram[16'h0ca2] = 8'hea; ram[16'h0ca3] = 8'hea; ram[16'h0ca4] = 8'h08; ram[16'h0ca5] = 8'hc9; ram[16'h0ca6] = 8'h68; ram[16'h0ca7] = 8'hd0; 
ram[16'h0ca8] = 8'hfe; ram[16'h0ca9] = 8'h68; ram[16'h0caa] = 8'h48; ram[16'h0cab] = 8'hc9; ram[16'h0cac] = 8'hff; ram[16'h0cad] = 8'hd0; ram[16'h0cae] = 8'hfe; ram[16'h0caf] = 8'h28; 
ram[16'h0cb0] = 8'hc0; ram[16'h0cb1] = 8'h42; ram[16'h0cb2] = 8'hd0; ram[16'h0cb3] = 8'hfe; ram[16'h0cb4] = 8'he0; ram[16'h0cb5] = 8'h00; ram[16'h0cb6] = 8'hd0; ram[16'h0cb7] = 8'hfe; 
ram[16'h0cb8] = 8'ha0; ram[16'h0cb9] = 8'h42; ram[16'h0cba] = 8'ha2; ram[16'h0cbb] = 8'h02; ram[16'h0cbc] = 8'h62; ram[16'h0cbd] = 8'hc8; ram[16'h0cbe] = 8'hca; ram[16'h0cbf] = 8'hca; 

ram[16'h0cc0] = 8'hd0; ram[16'h0cc1] = 8'hfe; ram[16'h0cc2] = 8'ha9; ram[16'h0cc3] = 8'h00; ram[16'h0cc4] = 8'h48; ram[16'h0cc5] = 8'ha9; ram[16'h0cc6] = 8'h9d; ram[16'h0cc7] = 8'h28; 
ram[16'h0cc8] = 8'h62; ram[16'h0cc9] = 8'hea; ram[16'h0cca] = 8'hea; ram[16'h0ccb] = 8'h08; ram[16'h0ccc] = 8'hc9; ram[16'h0ccd] = 8'h9d; ram[16'h0cce] = 8'hd0; ram[16'h0ccf] = 8'hfe; 
ram[16'h0cd0] = 8'h68; ram[16'h0cd1] = 8'h48; ram[16'h0cd2] = 8'hc9; ram[16'h0cd3] = 8'h30; ram[16'h0cd4] = 8'hd0; ram[16'h0cd5] = 8'hfe; ram[16'h0cd6] = 8'h28; ram[16'h0cd7] = 8'ha9; 
ram[16'h0cd8] = 8'hff; ram[16'h0cd9] = 8'h48; ram[16'h0cda] = 8'ha9; ram[16'h0cdb] = 8'h48; ram[16'h0cdc] = 8'h28; ram[16'h0cdd] = 8'h62; ram[16'h0cde] = 8'hea; ram[16'h0cdf] = 8'hea; 

ram[16'h0ce0] = 8'h08; ram[16'h0ce1] = 8'hc9; ram[16'h0ce2] = 8'h48; ram[16'h0ce3] = 8'hd0; ram[16'h0ce4] = 8'hfe; ram[16'h0ce5] = 8'h68; ram[16'h0ce6] = 8'h48; ram[16'h0ce7] = 8'hc9; 
ram[16'h0ce8] = 8'hff; ram[16'h0ce9] = 8'hd0; ram[16'h0cea] = 8'hfe; ram[16'h0ceb] = 8'h28; ram[16'h0cec] = 8'hc0; ram[16'h0ced] = 8'h42; ram[16'h0cee] = 8'hd0; ram[16'h0cef] = 8'hfe; 
ram[16'h0cf0] = 8'he0; ram[16'h0cf1] = 8'h00; ram[16'h0cf2] = 8'hd0; ram[16'h0cf3] = 8'hfe; ram[16'h0cf4] = 8'ha0; ram[16'h0cf5] = 8'h42; ram[16'h0cf6] = 8'ha2; ram[16'h0cf7] = 8'h02; 
ram[16'h0cf8] = 8'h82; ram[16'h0cf9] = 8'hc8; ram[16'h0cfa] = 8'hca; ram[16'h0cfb] = 8'hca; ram[16'h0cfc] = 8'hd0; ram[16'h0cfd] = 8'hfe; ram[16'h0cfe] = 8'ha9; ram[16'h0cff] = 8'h00; 

ram[16'h0d00] = 8'h48; ram[16'h0d01] = 8'ha9; ram[16'h0d02] = 8'h7d; ram[16'h0d03] = 8'h28; ram[16'h0d04] = 8'h82; ram[16'h0d05] = 8'hea; ram[16'h0d06] = 8'hea; ram[16'h0d07] = 8'h08; 
ram[16'h0d08] = 8'hc9; ram[16'h0d09] = 8'h7d; ram[16'h0d0a] = 8'hd0; ram[16'h0d0b] = 8'hfe; ram[16'h0d0c] = 8'h68; ram[16'h0d0d] = 8'h48; ram[16'h0d0e] = 8'hc9; ram[16'h0d0f] = 8'h30; 
ram[16'h0d10] = 8'hd0; ram[16'h0d11] = 8'hfe; ram[16'h0d12] = 8'h28; ram[16'h0d13] = 8'ha9; ram[16'h0d14] = 8'hff; ram[16'h0d15] = 8'h48; ram[16'h0d16] = 8'ha9; ram[16'h0d17] = 8'h28; 
ram[16'h0d18] = 8'h28; ram[16'h0d19] = 8'h82; ram[16'h0d1a] = 8'hea; ram[16'h0d1b] = 8'hea; ram[16'h0d1c] = 8'h08; ram[16'h0d1d] = 8'hc9; ram[16'h0d1e] = 8'h28; ram[16'h0d1f] = 8'hd0; 

ram[16'h0d20] = 8'hfe; ram[16'h0d21] = 8'h68; ram[16'h0d22] = 8'h48; ram[16'h0d23] = 8'hc9; ram[16'h0d24] = 8'hff; ram[16'h0d25] = 8'hd0; ram[16'h0d26] = 8'hfe; ram[16'h0d27] = 8'h28; 
ram[16'h0d28] = 8'hc0; ram[16'h0d29] = 8'h42; ram[16'h0d2a] = 8'hd0; ram[16'h0d2b] = 8'hfe; ram[16'h0d2c] = 8'he0; ram[16'h0d2d] = 8'h00; ram[16'h0d2e] = 8'hd0; ram[16'h0d2f] = 8'hfe; 
ram[16'h0d30] = 8'ha0; ram[16'h0d31] = 8'h42; ram[16'h0d32] = 8'ha2; ram[16'h0d33] = 8'h02; ram[16'h0d34] = 8'hc2; ram[16'h0d35] = 8'hc8; ram[16'h0d36] = 8'hca; ram[16'h0d37] = 8'hca; 
ram[16'h0d38] = 8'hd0; ram[16'h0d39] = 8'hfe; ram[16'h0d3a] = 8'ha9; ram[16'h0d3b] = 8'h00; ram[16'h0d3c] = 8'h48; ram[16'h0d3d] = 8'ha9; ram[16'h0d3e] = 8'h3d; ram[16'h0d3f] = 8'h28; 

ram[16'h0d40] = 8'hc2; ram[16'h0d41] = 8'hea; ram[16'h0d42] = 8'hea; ram[16'h0d43] = 8'h08; ram[16'h0d44] = 8'hc9; ram[16'h0d45] = 8'h3d; ram[16'h0d46] = 8'hd0; ram[16'h0d47] = 8'hfe; 
ram[16'h0d48] = 8'h68; ram[16'h0d49] = 8'h48; ram[16'h0d4a] = 8'hc9; ram[16'h0d4b] = 8'h30; ram[16'h0d4c] = 8'hd0; ram[16'h0d4d] = 8'hfe; ram[16'h0d4e] = 8'h28; ram[16'h0d4f] = 8'ha9; 
ram[16'h0d50] = 8'hff; ram[16'h0d51] = 8'h48; ram[16'h0d52] = 8'ha9; ram[16'h0d53] = 8'he8; ram[16'h0d54] = 8'h28; ram[16'h0d55] = 8'hc2; ram[16'h0d56] = 8'hea; ram[16'h0d57] = 8'hea; 
ram[16'h0d58] = 8'h08; ram[16'h0d59] = 8'hc9; ram[16'h0d5a] = 8'he8; ram[16'h0d5b] = 8'hd0; ram[16'h0d5c] = 8'hfe; ram[16'h0d5d] = 8'h68; ram[16'h0d5e] = 8'h48; ram[16'h0d5f] = 8'hc9; 

ram[16'h0d60] = 8'hff; ram[16'h0d61] = 8'hd0; ram[16'h0d62] = 8'hfe; ram[16'h0d63] = 8'h28; ram[16'h0d64] = 8'hc0; ram[16'h0d65] = 8'h42; ram[16'h0d66] = 8'hd0; ram[16'h0d67] = 8'hfe; 
ram[16'h0d68] = 8'he0; ram[16'h0d69] = 8'h00; ram[16'h0d6a] = 8'hd0; ram[16'h0d6b] = 8'hfe; ram[16'h0d6c] = 8'ha0; ram[16'h0d6d] = 8'h42; ram[16'h0d6e] = 8'ha2; ram[16'h0d6f] = 8'h02; 
ram[16'h0d70] = 8'he2; ram[16'h0d71] = 8'hc8; ram[16'h0d72] = 8'hca; ram[16'h0d73] = 8'hca; ram[16'h0d74] = 8'hd0; ram[16'h0d75] = 8'hfe; ram[16'h0d76] = 8'ha9; ram[16'h0d77] = 8'h00; 
ram[16'h0d78] = 8'h48; ram[16'h0d79] = 8'ha9; ram[16'h0d7a] = 8'h1d; ram[16'h0d7b] = 8'h28; ram[16'h0d7c] = 8'he2; ram[16'h0d7d] = 8'hea; ram[16'h0d7e] = 8'hea; ram[16'h0d7f] = 8'h08; 

ram[16'h0d80] = 8'hc9; ram[16'h0d81] = 8'h1d; ram[16'h0d82] = 8'hd0; ram[16'h0d83] = 8'hfe; ram[16'h0d84] = 8'h68; ram[16'h0d85] = 8'h48; ram[16'h0d86] = 8'hc9; ram[16'h0d87] = 8'h30; 
ram[16'h0d88] = 8'hd0; ram[16'h0d89] = 8'hfe; ram[16'h0d8a] = 8'h28; ram[16'h0d8b] = 8'ha9; ram[16'h0d8c] = 8'hff; ram[16'h0d8d] = 8'h48; ram[16'h0d8e] = 8'ha9; ram[16'h0d8f] = 8'hc8; 
ram[16'h0d90] = 8'h28; ram[16'h0d91] = 8'he2; ram[16'h0d92] = 8'hea; ram[16'h0d93] = 8'hea; ram[16'h0d94] = 8'h08; ram[16'h0d95] = 8'hc9; ram[16'h0d96] = 8'hc8; ram[16'h0d97] = 8'hd0; 
ram[16'h0d98] = 8'hfe; ram[16'h0d99] = 8'h68; ram[16'h0d9a] = 8'h48; ram[16'h0d9b] = 8'hc9; ram[16'h0d9c] = 8'hff; ram[16'h0d9d] = 8'hd0; ram[16'h0d9e] = 8'hfe; ram[16'h0d9f] = 8'h28; 

ram[16'h0da0] = 8'hc0; ram[16'h0da1] = 8'h42; ram[16'h0da2] = 8'hd0; ram[16'h0da3] = 8'hfe; ram[16'h0da4] = 8'he0; ram[16'h0da5] = 8'h00; ram[16'h0da6] = 8'hd0; ram[16'h0da7] = 8'hfe; 
ram[16'h0da8] = 8'ha0; ram[16'h0da9] = 8'h42; ram[16'h0daa] = 8'ha2; ram[16'h0dab] = 8'h02; ram[16'h0dac] = 8'h44; ram[16'h0dad] = 8'hc8; ram[16'h0dae] = 8'hca; ram[16'h0daf] = 8'hca; 
ram[16'h0db0] = 8'hd0; ram[16'h0db1] = 8'hfe; ram[16'h0db2] = 8'ha9; ram[16'h0db3] = 8'h00; ram[16'h0db4] = 8'h48; ram[16'h0db5] = 8'ha9; ram[16'h0db6] = 8'hbb; ram[16'h0db7] = 8'h28; 
ram[16'h0db8] = 8'h44; ram[16'h0db9] = 8'hea; ram[16'h0dba] = 8'hea; ram[16'h0dbb] = 8'h08; ram[16'h0dbc] = 8'hc9; ram[16'h0dbd] = 8'hbb; ram[16'h0dbe] = 8'hd0; ram[16'h0dbf] = 8'hfe; 

ram[16'h0dc0] = 8'h68; ram[16'h0dc1] = 8'h48; ram[16'h0dc2] = 8'hc9; ram[16'h0dc3] = 8'h30; ram[16'h0dc4] = 8'hd0; ram[16'h0dc5] = 8'hfe; ram[16'h0dc6] = 8'h28; ram[16'h0dc7] = 8'ha9; 
ram[16'h0dc8] = 8'hff; ram[16'h0dc9] = 8'h48; ram[16'h0dca] = 8'ha9; ram[16'h0dcb] = 8'h66; ram[16'h0dcc] = 8'h28; ram[16'h0dcd] = 8'h44; ram[16'h0dce] = 8'hea; ram[16'h0dcf] = 8'hea; 
ram[16'h0dd0] = 8'h08; ram[16'h0dd1] = 8'hc9; ram[16'h0dd2] = 8'h66; ram[16'h0dd3] = 8'hd0; ram[16'h0dd4] = 8'hfe; ram[16'h0dd5] = 8'h68; ram[16'h0dd6] = 8'h48; ram[16'h0dd7] = 8'hc9; 
ram[16'h0dd8] = 8'hff; ram[16'h0dd9] = 8'hd0; ram[16'h0dda] = 8'hfe; ram[16'h0ddb] = 8'h28; ram[16'h0ddc] = 8'hc0; ram[16'h0ddd] = 8'h42; ram[16'h0dde] = 8'hd0; ram[16'h0ddf] = 8'hfe; 

ram[16'h0de0] = 8'he0; ram[16'h0de1] = 8'h00; ram[16'h0de2] = 8'hd0; ram[16'h0de3] = 8'hfe; ram[16'h0de4] = 8'ha0; ram[16'h0de5] = 8'h42; ram[16'h0de6] = 8'ha2; ram[16'h0de7] = 8'h02; 
ram[16'h0de8] = 8'h54; ram[16'h0de9] = 8'hc8; ram[16'h0dea] = 8'hca; ram[16'h0deb] = 8'hca; ram[16'h0dec] = 8'hd0; ram[16'h0ded] = 8'hfe; ram[16'h0dee] = 8'ha9; ram[16'h0def] = 8'h00; 
ram[16'h0df0] = 8'h48; ram[16'h0df1] = 8'ha9; ram[16'h0df2] = 8'hab; ram[16'h0df3] = 8'h28; ram[16'h0df4] = 8'h54; ram[16'h0df5] = 8'hea; ram[16'h0df6] = 8'hea; ram[16'h0df7] = 8'h08; 
ram[16'h0df8] = 8'hc9; ram[16'h0df9] = 8'hab; ram[16'h0dfa] = 8'hd0; ram[16'h0dfb] = 8'hfe; ram[16'h0dfc] = 8'h68; ram[16'h0dfd] = 8'h48; ram[16'h0dfe] = 8'hc9; ram[16'h0dff] = 8'h30; 

ram[16'h0e00] = 8'hd0; ram[16'h0e01] = 8'hfe; ram[16'h0e02] = 8'h28; ram[16'h0e03] = 8'ha9; ram[16'h0e04] = 8'hff; ram[16'h0e05] = 8'h48; ram[16'h0e06] = 8'ha9; ram[16'h0e07] = 8'h56; 
ram[16'h0e08] = 8'h28; ram[16'h0e09] = 8'h54; ram[16'h0e0a] = 8'hea; ram[16'h0e0b] = 8'hea; ram[16'h0e0c] = 8'h08; ram[16'h0e0d] = 8'hc9; ram[16'h0e0e] = 8'h56; ram[16'h0e0f] = 8'hd0; 
ram[16'h0e10] = 8'hfe; ram[16'h0e11] = 8'h68; ram[16'h0e12] = 8'h48; ram[16'h0e13] = 8'hc9; ram[16'h0e14] = 8'hff; ram[16'h0e15] = 8'hd0; ram[16'h0e16] = 8'hfe; ram[16'h0e17] = 8'h28; 
ram[16'h0e18] = 8'hc0; ram[16'h0e19] = 8'h42; ram[16'h0e1a] = 8'hd0; ram[16'h0e1b] = 8'hfe; ram[16'h0e1c] = 8'he0; ram[16'h0e1d] = 8'h00; ram[16'h0e1e] = 8'hd0; ram[16'h0e1f] = 8'hfe; 

ram[16'h0e20] = 8'ha0; ram[16'h0e21] = 8'h42; ram[16'h0e22] = 8'ha2; ram[16'h0e23] = 8'h02; ram[16'h0e24] = 8'hd4; ram[16'h0e25] = 8'hc8; ram[16'h0e26] = 8'hca; ram[16'h0e27] = 8'hca; 
ram[16'h0e28] = 8'hd0; ram[16'h0e29] = 8'hfe; ram[16'h0e2a] = 8'ha9; ram[16'h0e2b] = 8'h00; ram[16'h0e2c] = 8'h48; ram[16'h0e2d] = 8'ha9; ram[16'h0e2e] = 8'h2b; ram[16'h0e2f] = 8'h28; 
ram[16'h0e30] = 8'hd4; ram[16'h0e31] = 8'hea; ram[16'h0e32] = 8'hea; ram[16'h0e33] = 8'h08; ram[16'h0e34] = 8'hc9; ram[16'h0e35] = 8'h2b; ram[16'h0e36] = 8'hd0; ram[16'h0e37] = 8'hfe; 
ram[16'h0e38] = 8'h68; ram[16'h0e39] = 8'h48; ram[16'h0e3a] = 8'hc9; ram[16'h0e3b] = 8'h30; ram[16'h0e3c] = 8'hd0; ram[16'h0e3d] = 8'hfe; ram[16'h0e3e] = 8'h28; ram[16'h0e3f] = 8'ha9; 

ram[16'h0e40] = 8'hff; ram[16'h0e41] = 8'h48; ram[16'h0e42] = 8'ha9; ram[16'h0e43] = 8'hd6; ram[16'h0e44] = 8'h28; ram[16'h0e45] = 8'hd4; ram[16'h0e46] = 8'hea; ram[16'h0e47] = 8'hea; 
ram[16'h0e48] = 8'h08; ram[16'h0e49] = 8'hc9; ram[16'h0e4a] = 8'hd6; ram[16'h0e4b] = 8'hd0; ram[16'h0e4c] = 8'hfe; ram[16'h0e4d] = 8'h68; ram[16'h0e4e] = 8'h48; ram[16'h0e4f] = 8'hc9; 
ram[16'h0e50] = 8'hff; ram[16'h0e51] = 8'hd0; ram[16'h0e52] = 8'hfe; ram[16'h0e53] = 8'h28; ram[16'h0e54] = 8'hc0; ram[16'h0e55] = 8'h42; ram[16'h0e56] = 8'hd0; ram[16'h0e57] = 8'hfe; 
ram[16'h0e58] = 8'he0; ram[16'h0e59] = 8'h00; ram[16'h0e5a] = 8'hd0; ram[16'h0e5b] = 8'hfe; ram[16'h0e5c] = 8'ha0; ram[16'h0e5d] = 8'h42; ram[16'h0e5e] = 8'ha2; ram[16'h0e5f] = 8'h02; 

ram[16'h0e60] = 8'hf4; ram[16'h0e61] = 8'hc8; ram[16'h0e62] = 8'hca; ram[16'h0e63] = 8'hca; ram[16'h0e64] = 8'hd0; ram[16'h0e65] = 8'hfe; ram[16'h0e66] = 8'ha9; ram[16'h0e67] = 8'h00; 
ram[16'h0e68] = 8'h48; ram[16'h0e69] = 8'ha9; ram[16'h0e6a] = 8'h0b; ram[16'h0e6b] = 8'h28; ram[16'h0e6c] = 8'hf4; ram[16'h0e6d] = 8'hea; ram[16'h0e6e] = 8'hea; ram[16'h0e6f] = 8'h08; 
ram[16'h0e70] = 8'hc9; ram[16'h0e71] = 8'h0b; ram[16'h0e72] = 8'hd0; ram[16'h0e73] = 8'hfe; ram[16'h0e74] = 8'h68; ram[16'h0e75] = 8'h48; ram[16'h0e76] = 8'hc9; ram[16'h0e77] = 8'h30; 
ram[16'h0e78] = 8'hd0; ram[16'h0e79] = 8'hfe; ram[16'h0e7a] = 8'h28; ram[16'h0e7b] = 8'ha9; ram[16'h0e7c] = 8'hff; ram[16'h0e7d] = 8'h48; ram[16'h0e7e] = 8'ha9; ram[16'h0e7f] = 8'hb6; 

ram[16'h0e80] = 8'h28; ram[16'h0e81] = 8'hf4; ram[16'h0e82] = 8'hea; ram[16'h0e83] = 8'hea; ram[16'h0e84] = 8'h08; ram[16'h0e85] = 8'hc9; ram[16'h0e86] = 8'hb6; ram[16'h0e87] = 8'hd0; 
ram[16'h0e88] = 8'hfe; ram[16'h0e89] = 8'h68; ram[16'h0e8a] = 8'h48; ram[16'h0e8b] = 8'hc9; ram[16'h0e8c] = 8'hff; ram[16'h0e8d] = 8'hd0; ram[16'h0e8e] = 8'hfe; ram[16'h0e8f] = 8'h28; 
ram[16'h0e90] = 8'hc0; ram[16'h0e91] = 8'h42; ram[16'h0e92] = 8'hd0; ram[16'h0e93] = 8'hfe; ram[16'h0e94] = 8'he0; ram[16'h0e95] = 8'h00; ram[16'h0e96] = 8'hd0; ram[16'h0e97] = 8'hfe; 
ram[16'h0e98] = 8'ha0; ram[16'h0e99] = 8'h42; ram[16'h0e9a] = 8'ha2; ram[16'h0e9b] = 8'h01; ram[16'h0e9c] = 8'h5c; ram[16'h0e9d] = 8'hc8; ram[16'h0e9e] = 8'hc8; ram[16'h0e9f] = 8'hca; 

ram[16'h0ea0] = 8'hd0; ram[16'h0ea1] = 8'hfe; ram[16'h0ea2] = 8'ha9; ram[16'h0ea3] = 8'h00; ram[16'h0ea4] = 8'h48; ram[16'h0ea5] = 8'ha9; ram[16'h0ea6] = 8'ha3; ram[16'h0ea7] = 8'h28; 
ram[16'h0ea8] = 8'h5c; ram[16'h0ea9] = 8'hea; ram[16'h0eaa] = 8'hea; ram[16'h0eab] = 8'h08; ram[16'h0eac] = 8'hc9; ram[16'h0ead] = 8'ha3; ram[16'h0eae] = 8'hd0; ram[16'h0eaf] = 8'hfe; 
ram[16'h0eb0] = 8'h68; ram[16'h0eb1] = 8'h48; ram[16'h0eb2] = 8'hc9; ram[16'h0eb3] = 8'h30; ram[16'h0eb4] = 8'hd0; ram[16'h0eb5] = 8'hfe; ram[16'h0eb6] = 8'h28; ram[16'h0eb7] = 8'ha9; 
ram[16'h0eb8] = 8'hff; ram[16'h0eb9] = 8'h48; ram[16'h0eba] = 8'ha9; ram[16'h0ebb] = 8'h4e; ram[16'h0ebc] = 8'h28; ram[16'h0ebd] = 8'h5c; ram[16'h0ebe] = 8'hea; ram[16'h0ebf] = 8'hea; 

ram[16'h0ec0] = 8'h08; ram[16'h0ec1] = 8'hc9; ram[16'h0ec2] = 8'h4e; ram[16'h0ec3] = 8'hd0; ram[16'h0ec4] = 8'hfe; ram[16'h0ec5] = 8'h68; ram[16'h0ec6] = 8'h48; ram[16'h0ec7] = 8'hc9; 
ram[16'h0ec8] = 8'hff; ram[16'h0ec9] = 8'hd0; ram[16'h0eca] = 8'hfe; ram[16'h0ecb] = 8'h28; ram[16'h0ecc] = 8'hc0; ram[16'h0ecd] = 8'h42; ram[16'h0ece] = 8'hd0; ram[16'h0ecf] = 8'hfe; 
ram[16'h0ed0] = 8'he0; ram[16'h0ed1] = 8'h00; ram[16'h0ed2] = 8'hd0; ram[16'h0ed3] = 8'hfe; ram[16'h0ed4] = 8'ha0; ram[16'h0ed5] = 8'h42; ram[16'h0ed6] = 8'ha2; ram[16'h0ed7] = 8'h01; 
ram[16'h0ed8] = 8'hdc; ram[16'h0ed9] = 8'hc8; ram[16'h0eda] = 8'hc8; ram[16'h0edb] = 8'hca; ram[16'h0edc] = 8'hd0; ram[16'h0edd] = 8'hfe; ram[16'h0ede] = 8'ha9; ram[16'h0edf] = 8'h00; 

ram[16'h0ee0] = 8'h48; ram[16'h0ee1] = 8'ha9; ram[16'h0ee2] = 8'h23; ram[16'h0ee3] = 8'h28; ram[16'h0ee4] = 8'hdc; ram[16'h0ee5] = 8'hea; ram[16'h0ee6] = 8'hea; ram[16'h0ee7] = 8'h08; 
ram[16'h0ee8] = 8'hc9; ram[16'h0ee9] = 8'h23; ram[16'h0eea] = 8'hd0; ram[16'h0eeb] = 8'hfe; ram[16'h0eec] = 8'h68; ram[16'h0eed] = 8'h48; ram[16'h0eee] = 8'hc9; ram[16'h0eef] = 8'h30; 
ram[16'h0ef0] = 8'hd0; ram[16'h0ef1] = 8'hfe; ram[16'h0ef2] = 8'h28; ram[16'h0ef3] = 8'ha9; ram[16'h0ef4] = 8'hff; ram[16'h0ef5] = 8'h48; ram[16'h0ef6] = 8'ha9; ram[16'h0ef7] = 8'hce; 
ram[16'h0ef8] = 8'h28; ram[16'h0ef9] = 8'hdc; ram[16'h0efa] = 8'hea; ram[16'h0efb] = 8'hea; ram[16'h0efc] = 8'h08; ram[16'h0efd] = 8'hc9; ram[16'h0efe] = 8'hce; ram[16'h0eff] = 8'hd0; 

ram[16'h0f00] = 8'hfe; ram[16'h0f01] = 8'h68; ram[16'h0f02] = 8'h48; ram[16'h0f03] = 8'hc9; ram[16'h0f04] = 8'hff; ram[16'h0f05] = 8'hd0; ram[16'h0f06] = 8'hfe; ram[16'h0f07] = 8'h28; 
ram[16'h0f08] = 8'hc0; ram[16'h0f09] = 8'h42; ram[16'h0f0a] = 8'hd0; ram[16'h0f0b] = 8'hfe; ram[16'h0f0c] = 8'he0; ram[16'h0f0d] = 8'h00; ram[16'h0f0e] = 8'hd0; ram[16'h0f0f] = 8'hfe; 
ram[16'h0f10] = 8'ha0; ram[16'h0f11] = 8'h42; ram[16'h0f12] = 8'ha2; ram[16'h0f13] = 8'h01; ram[16'h0f14] = 8'hfc; ram[16'h0f15] = 8'hc8; ram[16'h0f16] = 8'hc8; ram[16'h0f17] = 8'hca; 
ram[16'h0f18] = 8'hd0; ram[16'h0f19] = 8'hfe; ram[16'h0f1a] = 8'ha9; ram[16'h0f1b] = 8'h00; ram[16'h0f1c] = 8'h48; ram[16'h0f1d] = 8'ha9; ram[16'h0f1e] = 8'h03; ram[16'h0f1f] = 8'h28; 

ram[16'h0f20] = 8'hfc; ram[16'h0f21] = 8'hea; ram[16'h0f22] = 8'hea; ram[16'h0f23] = 8'h08; ram[16'h0f24] = 8'hc9; ram[16'h0f25] = 8'h03; ram[16'h0f26] = 8'hd0; ram[16'h0f27] = 8'hfe; 
ram[16'h0f28] = 8'h68; ram[16'h0f29] = 8'h48; ram[16'h0f2a] = 8'hc9; ram[16'h0f2b] = 8'h30; ram[16'h0f2c] = 8'hd0; ram[16'h0f2d] = 8'hfe; ram[16'h0f2e] = 8'h28; ram[16'h0f2f] = 8'ha9; 
ram[16'h0f30] = 8'hff; ram[16'h0f31] = 8'h48; ram[16'h0f32] = 8'ha9; ram[16'h0f33] = 8'hae; ram[16'h0f34] = 8'h28; ram[16'h0f35] = 8'hfc; ram[16'h0f36] = 8'hea; ram[16'h0f37] = 8'hea; 
ram[16'h0f38] = 8'h08; ram[16'h0f39] = 8'hc9; ram[16'h0f3a] = 8'hae; ram[16'h0f3b] = 8'hd0; ram[16'h0f3c] = 8'hfe; ram[16'h0f3d] = 8'h68; ram[16'h0f3e] = 8'h48; ram[16'h0f3f] = 8'hc9; 

ram[16'h0f40] = 8'hff; ram[16'h0f41] = 8'hd0; ram[16'h0f42] = 8'hfe; ram[16'h0f43] = 8'h28; ram[16'h0f44] = 8'hc0; ram[16'h0f45] = 8'h42; ram[16'h0f46] = 8'hd0; ram[16'h0f47] = 8'hfe; 
ram[16'h0f48] = 8'he0; ram[16'h0f49] = 8'h00; ram[16'h0f4a] = 8'hd0; ram[16'h0f4b] = 8'hfe; ram[16'h0f4c] = 8'ha0; ram[16'h0f4d] = 8'h42; ram[16'h0f4e] = 8'ha2; ram[16'h0f4f] = 8'h03; 
ram[16'h0f50] = 8'h03; ram[16'h0f51] = 8'hca; ram[16'h0f52] = 8'hca; ram[16'h0f53] = 8'hca; ram[16'h0f54] = 8'hd0; ram[16'h0f55] = 8'hfe; ram[16'h0f56] = 8'ha9; ram[16'h0f57] = 8'h00; 
ram[16'h0f58] = 8'h48; ram[16'h0f59] = 8'ha9; ram[16'h0f5a] = 8'hfc; ram[16'h0f5b] = 8'h28; ram[16'h0f5c] = 8'h03; ram[16'h0f5d] = 8'hea; ram[16'h0f5e] = 8'hea; ram[16'h0f5f] = 8'h08; 

ram[16'h0f60] = 8'hc9; ram[16'h0f61] = 8'hfc; ram[16'h0f62] = 8'hd0; ram[16'h0f63] = 8'hfe; ram[16'h0f64] = 8'h68; ram[16'h0f65] = 8'h48; ram[16'h0f66] = 8'hc9; ram[16'h0f67] = 8'h30; 
ram[16'h0f68] = 8'hd0; ram[16'h0f69] = 8'hfe; ram[16'h0f6a] = 8'h28; ram[16'h0f6b] = 8'ha9; ram[16'h0f6c] = 8'hff; ram[16'h0f6d] = 8'h48; ram[16'h0f6e] = 8'ha9; ram[16'h0f6f] = 8'ha7; 
ram[16'h0f70] = 8'h28; ram[16'h0f71] = 8'h03; ram[16'h0f72] = 8'hea; ram[16'h0f73] = 8'hea; ram[16'h0f74] = 8'h08; ram[16'h0f75] = 8'hc9; ram[16'h0f76] = 8'ha7; ram[16'h0f77] = 8'hd0; 
ram[16'h0f78] = 8'hfe; ram[16'h0f79] = 8'h68; ram[16'h0f7a] = 8'h48; ram[16'h0f7b] = 8'hc9; ram[16'h0f7c] = 8'hff; ram[16'h0f7d] = 8'hd0; ram[16'h0f7e] = 8'hfe; ram[16'h0f7f] = 8'h28; 

ram[16'h0f80] = 8'hc0; ram[16'h0f81] = 8'h42; ram[16'h0f82] = 8'hd0; ram[16'h0f83] = 8'hfe; ram[16'h0f84] = 8'he0; ram[16'h0f85] = 8'h00; ram[16'h0f86] = 8'hd0; ram[16'h0f87] = 8'hfe; 
ram[16'h0f88] = 8'ha0; ram[16'h0f89] = 8'h42; ram[16'h0f8a] = 8'ha2; ram[16'h0f8b] = 8'h03; ram[16'h0f8c] = 8'h13; ram[16'h0f8d] = 8'hca; ram[16'h0f8e] = 8'hca; ram[16'h0f8f] = 8'hca; 
ram[16'h0f90] = 8'hd0; ram[16'h0f91] = 8'hfe; ram[16'h0f92] = 8'ha9; ram[16'h0f93] = 8'h00; ram[16'h0f94] = 8'h48; ram[16'h0f95] = 8'ha9; ram[16'h0f96] = 8'hec; ram[16'h0f97] = 8'h28; 
ram[16'h0f98] = 8'h13; ram[16'h0f99] = 8'hea; ram[16'h0f9a] = 8'hea; ram[16'h0f9b] = 8'h08; ram[16'h0f9c] = 8'hc9; ram[16'h0f9d] = 8'hec; ram[16'h0f9e] = 8'hd0; ram[16'h0f9f] = 8'hfe; 

ram[16'h0fa0] = 8'h68; ram[16'h0fa1] = 8'h48; ram[16'h0fa2] = 8'hc9; ram[16'h0fa3] = 8'h30; ram[16'h0fa4] = 8'hd0; ram[16'h0fa5] = 8'hfe; ram[16'h0fa6] = 8'h28; ram[16'h0fa7] = 8'ha9; 
ram[16'h0fa8] = 8'hff; ram[16'h0fa9] = 8'h48; ram[16'h0faa] = 8'ha9; ram[16'h0fab] = 8'h97; ram[16'h0fac] = 8'h28; ram[16'h0fad] = 8'h13; ram[16'h0fae] = 8'hea; ram[16'h0faf] = 8'hea; 
ram[16'h0fb0] = 8'h08; ram[16'h0fb1] = 8'hc9; ram[16'h0fb2] = 8'h97; ram[16'h0fb3] = 8'hd0; ram[16'h0fb4] = 8'hfe; ram[16'h0fb5] = 8'h68; ram[16'h0fb6] = 8'h48; ram[16'h0fb7] = 8'hc9; 
ram[16'h0fb8] = 8'hff; ram[16'h0fb9] = 8'hd0; ram[16'h0fba] = 8'hfe; ram[16'h0fbb] = 8'h28; ram[16'h0fbc] = 8'hc0; ram[16'h0fbd] = 8'h42; ram[16'h0fbe] = 8'hd0; ram[16'h0fbf] = 8'hfe; 

ram[16'h0fc0] = 8'he0; ram[16'h0fc1] = 8'h00; ram[16'h0fc2] = 8'hd0; ram[16'h0fc3] = 8'hfe; ram[16'h0fc4] = 8'ha0; ram[16'h0fc5] = 8'h42; ram[16'h0fc6] = 8'ha2; ram[16'h0fc7] = 8'h03; 
ram[16'h0fc8] = 8'h23; ram[16'h0fc9] = 8'hca; ram[16'h0fca] = 8'hca; ram[16'h0fcb] = 8'hca; ram[16'h0fcc] = 8'hd0; ram[16'h0fcd] = 8'hfe; ram[16'h0fce] = 8'ha9; ram[16'h0fcf] = 8'h00; 
ram[16'h0fd0] = 8'h48; ram[16'h0fd1] = 8'ha9; ram[16'h0fd2] = 8'hdc; ram[16'h0fd3] = 8'h28; ram[16'h0fd4] = 8'h23; ram[16'h0fd5] = 8'hea; ram[16'h0fd6] = 8'hea; ram[16'h0fd7] = 8'h08; 
ram[16'h0fd8] = 8'hc9; ram[16'h0fd9] = 8'hdc; ram[16'h0fda] = 8'hd0; ram[16'h0fdb] = 8'hfe; ram[16'h0fdc] = 8'h68; ram[16'h0fdd] = 8'h48; ram[16'h0fde] = 8'hc9; ram[16'h0fdf] = 8'h30; 

ram[16'h0fe0] = 8'hd0; ram[16'h0fe1] = 8'hfe; ram[16'h0fe2] = 8'h28; ram[16'h0fe3] = 8'ha9; ram[16'h0fe4] = 8'hff; ram[16'h0fe5] = 8'h48; ram[16'h0fe6] = 8'ha9; ram[16'h0fe7] = 8'h87; 
ram[16'h0fe8] = 8'h28; ram[16'h0fe9] = 8'h23; ram[16'h0fea] = 8'hea; ram[16'h0feb] = 8'hea; ram[16'h0fec] = 8'h08; ram[16'h0fed] = 8'hc9; ram[16'h0fee] = 8'h87; ram[16'h0fef] = 8'hd0; 
ram[16'h0ff0] = 8'hfe; ram[16'h0ff1] = 8'h68; ram[16'h0ff2] = 8'h48; ram[16'h0ff3] = 8'hc9; ram[16'h0ff4] = 8'hff; ram[16'h0ff5] = 8'hd0; ram[16'h0ff6] = 8'hfe; ram[16'h0ff7] = 8'h28; 
ram[16'h0ff8] = 8'hc0; ram[16'h0ff9] = 8'h42; ram[16'h0ffa] = 8'hd0; ram[16'h0ffb] = 8'hfe; ram[16'h0ffc] = 8'he0; ram[16'h0ffd] = 8'h00; ram[16'h0ffe] = 8'hd0; ram[16'h0fff] = 8'hfe; 

ram[16'h1000] = 8'ha0; ram[16'h1001] = 8'h42; ram[16'h1002] = 8'ha2; ram[16'h1003] = 8'h03; ram[16'h1004] = 8'h33; ram[16'h1005] = 8'hca; ram[16'h1006] = 8'hca; ram[16'h1007] = 8'hca; 
ram[16'h1008] = 8'hd0; ram[16'h1009] = 8'hfe; ram[16'h100a] = 8'ha9; ram[16'h100b] = 8'h00; ram[16'h100c] = 8'h48; ram[16'h100d] = 8'ha9; ram[16'h100e] = 8'hcc; ram[16'h100f] = 8'h28; 
ram[16'h1010] = 8'h33; ram[16'h1011] = 8'hea; ram[16'h1012] = 8'hea; ram[16'h1013] = 8'h08; ram[16'h1014] = 8'hc9; ram[16'h1015] = 8'hcc; ram[16'h1016] = 8'hd0; ram[16'h1017] = 8'hfe; 
ram[16'h1018] = 8'h68; ram[16'h1019] = 8'h48; ram[16'h101a] = 8'hc9; ram[16'h101b] = 8'h30; ram[16'h101c] = 8'hd0; ram[16'h101d] = 8'hfe; ram[16'h101e] = 8'h28; ram[16'h101f] = 8'ha9; 

ram[16'h1020] = 8'hff; ram[16'h1021] = 8'h48; ram[16'h1022] = 8'ha9; ram[16'h1023] = 8'h77; ram[16'h1024] = 8'h28; ram[16'h1025] = 8'h33; ram[16'h1026] = 8'hea; ram[16'h1027] = 8'hea; 
ram[16'h1028] = 8'h08; ram[16'h1029] = 8'hc9; ram[16'h102a] = 8'h77; ram[16'h102b] = 8'hd0; ram[16'h102c] = 8'hfe; ram[16'h102d] = 8'h68; ram[16'h102e] = 8'h48; ram[16'h102f] = 8'hc9; 
ram[16'h1030] = 8'hff; ram[16'h1031] = 8'hd0; ram[16'h1032] = 8'hfe; ram[16'h1033] = 8'h28; ram[16'h1034] = 8'hc0; ram[16'h1035] = 8'h42; ram[16'h1036] = 8'hd0; ram[16'h1037] = 8'hfe; 
ram[16'h1038] = 8'he0; ram[16'h1039] = 8'h00; ram[16'h103a] = 8'hd0; ram[16'h103b] = 8'hfe; ram[16'h103c] = 8'ha0; ram[16'h103d] = 8'h42; ram[16'h103e] = 8'ha2; ram[16'h103f] = 8'h03; 

ram[16'h1040] = 8'h43; ram[16'h1041] = 8'hca; ram[16'h1042] = 8'hca; ram[16'h1043] = 8'hca; ram[16'h1044] = 8'hd0; ram[16'h1045] = 8'hfe; ram[16'h1046] = 8'ha9; ram[16'h1047] = 8'h00; 
ram[16'h1048] = 8'h48; ram[16'h1049] = 8'ha9; ram[16'h104a] = 8'hbc; ram[16'h104b] = 8'h28; ram[16'h104c] = 8'h43; ram[16'h104d] = 8'hea; ram[16'h104e] = 8'hea; ram[16'h104f] = 8'h08; 
ram[16'h1050] = 8'hc9; ram[16'h1051] = 8'hbc; ram[16'h1052] = 8'hd0; ram[16'h1053] = 8'hfe; ram[16'h1054] = 8'h68; ram[16'h1055] = 8'h48; ram[16'h1056] = 8'hc9; ram[16'h1057] = 8'h30; 
ram[16'h1058] = 8'hd0; ram[16'h1059] = 8'hfe; ram[16'h105a] = 8'h28; ram[16'h105b] = 8'ha9; ram[16'h105c] = 8'hff; ram[16'h105d] = 8'h48; ram[16'h105e] = 8'ha9; ram[16'h105f] = 8'h67; 

ram[16'h1060] = 8'h28; ram[16'h1061] = 8'h43; ram[16'h1062] = 8'hea; ram[16'h1063] = 8'hea; ram[16'h1064] = 8'h08; ram[16'h1065] = 8'hc9; ram[16'h1066] = 8'h67; ram[16'h1067] = 8'hd0; 
ram[16'h1068] = 8'hfe; ram[16'h1069] = 8'h68; ram[16'h106a] = 8'h48; ram[16'h106b] = 8'hc9; ram[16'h106c] = 8'hff; ram[16'h106d] = 8'hd0; ram[16'h106e] = 8'hfe; ram[16'h106f] = 8'h28; 
ram[16'h1070] = 8'hc0; ram[16'h1071] = 8'h42; ram[16'h1072] = 8'hd0; ram[16'h1073] = 8'hfe; ram[16'h1074] = 8'he0; ram[16'h1075] = 8'h00; ram[16'h1076] = 8'hd0; ram[16'h1077] = 8'hfe; 
ram[16'h1078] = 8'ha0; ram[16'h1079] = 8'h42; ram[16'h107a] = 8'ha2; ram[16'h107b] = 8'h03; ram[16'h107c] = 8'h53; ram[16'h107d] = 8'hca; ram[16'h107e] = 8'hca; ram[16'h107f] = 8'hca; 

ram[16'h1080] = 8'hd0; ram[16'h1081] = 8'hfe; ram[16'h1082] = 8'ha9; ram[16'h1083] = 8'h00; ram[16'h1084] = 8'h48; ram[16'h1085] = 8'ha9; ram[16'h1086] = 8'hac; ram[16'h1087] = 8'h28; 
ram[16'h1088] = 8'h53; ram[16'h1089] = 8'hea; ram[16'h108a] = 8'hea; ram[16'h108b] = 8'h08; ram[16'h108c] = 8'hc9; ram[16'h108d] = 8'hac; ram[16'h108e] = 8'hd0; ram[16'h108f] = 8'hfe; 
ram[16'h1090] = 8'h68; ram[16'h1091] = 8'h48; ram[16'h1092] = 8'hc9; ram[16'h1093] = 8'h30; ram[16'h1094] = 8'hd0; ram[16'h1095] = 8'hfe; ram[16'h1096] = 8'h28; ram[16'h1097] = 8'ha9; 
ram[16'h1098] = 8'hff; ram[16'h1099] = 8'h48; ram[16'h109a] = 8'ha9; ram[16'h109b] = 8'h57; ram[16'h109c] = 8'h28; ram[16'h109d] = 8'h53; ram[16'h109e] = 8'hea; ram[16'h109f] = 8'hea; 

ram[16'h10a0] = 8'h08; ram[16'h10a1] = 8'hc9; ram[16'h10a2] = 8'h57; ram[16'h10a3] = 8'hd0; ram[16'h10a4] = 8'hfe; ram[16'h10a5] = 8'h68; ram[16'h10a6] = 8'h48; ram[16'h10a7] = 8'hc9; 
ram[16'h10a8] = 8'hff; ram[16'h10a9] = 8'hd0; ram[16'h10aa] = 8'hfe; ram[16'h10ab] = 8'h28; ram[16'h10ac] = 8'hc0; ram[16'h10ad] = 8'h42; ram[16'h10ae] = 8'hd0; ram[16'h10af] = 8'hfe; 
ram[16'h10b0] = 8'he0; ram[16'h10b1] = 8'h00; ram[16'h10b2] = 8'hd0; ram[16'h10b3] = 8'hfe; ram[16'h10b4] = 8'ha0; ram[16'h10b5] = 8'h42; ram[16'h10b6] = 8'ha2; ram[16'h10b7] = 8'h03; 
ram[16'h10b8] = 8'h63; ram[16'h10b9] = 8'hca; ram[16'h10ba] = 8'hca; ram[16'h10bb] = 8'hca; ram[16'h10bc] = 8'hd0; ram[16'h10bd] = 8'hfe; ram[16'h10be] = 8'ha9; ram[16'h10bf] = 8'h00; 

ram[16'h10c0] = 8'h48; ram[16'h10c1] = 8'ha9; ram[16'h10c2] = 8'h9c; ram[16'h10c3] = 8'h28; ram[16'h10c4] = 8'h63; ram[16'h10c5] = 8'hea; ram[16'h10c6] = 8'hea; ram[16'h10c7] = 8'h08; 
ram[16'h10c8] = 8'hc9; ram[16'h10c9] = 8'h9c; ram[16'h10ca] = 8'hd0; ram[16'h10cb] = 8'hfe; ram[16'h10cc] = 8'h68; ram[16'h10cd] = 8'h48; ram[16'h10ce] = 8'hc9; ram[16'h10cf] = 8'h30; 
ram[16'h10d0] = 8'hd0; ram[16'h10d1] = 8'hfe; ram[16'h10d2] = 8'h28; ram[16'h10d3] = 8'ha9; ram[16'h10d4] = 8'hff; ram[16'h10d5] = 8'h48; ram[16'h10d6] = 8'ha9; ram[16'h10d7] = 8'h47; 
ram[16'h10d8] = 8'h28; ram[16'h10d9] = 8'h63; ram[16'h10da] = 8'hea; ram[16'h10db] = 8'hea; ram[16'h10dc] = 8'h08; ram[16'h10dd] = 8'hc9; ram[16'h10de] = 8'h47; ram[16'h10df] = 8'hd0; 

ram[16'h10e0] = 8'hfe; ram[16'h10e1] = 8'h68; ram[16'h10e2] = 8'h48; ram[16'h10e3] = 8'hc9; ram[16'h10e4] = 8'hff; ram[16'h10e5] = 8'hd0; ram[16'h10e6] = 8'hfe; ram[16'h10e7] = 8'h28; 
ram[16'h10e8] = 8'hc0; ram[16'h10e9] = 8'h42; ram[16'h10ea] = 8'hd0; ram[16'h10eb] = 8'hfe; ram[16'h10ec] = 8'he0; ram[16'h10ed] = 8'h00; ram[16'h10ee] = 8'hd0; ram[16'h10ef] = 8'hfe; 
ram[16'h10f0] = 8'ha0; ram[16'h10f1] = 8'h42; ram[16'h10f2] = 8'ha2; ram[16'h10f3] = 8'h03; ram[16'h10f4] = 8'h73; ram[16'h10f5] = 8'hca; ram[16'h10f6] = 8'hca; ram[16'h10f7] = 8'hca; 
ram[16'h10f8] = 8'hd0; ram[16'h10f9] = 8'hfe; ram[16'h10fa] = 8'ha9; ram[16'h10fb] = 8'h00; ram[16'h10fc] = 8'h48; ram[16'h10fd] = 8'ha9; ram[16'h10fe] = 8'h8c; ram[16'h10ff] = 8'h28; 

ram[16'h1100] = 8'h73; ram[16'h1101] = 8'hea; ram[16'h1102] = 8'hea; ram[16'h1103] = 8'h08; ram[16'h1104] = 8'hc9; ram[16'h1105] = 8'h8c; ram[16'h1106] = 8'hd0; ram[16'h1107] = 8'hfe; 
ram[16'h1108] = 8'h68; ram[16'h1109] = 8'h48; ram[16'h110a] = 8'hc9; ram[16'h110b] = 8'h30; ram[16'h110c] = 8'hd0; ram[16'h110d] = 8'hfe; ram[16'h110e] = 8'h28; ram[16'h110f] = 8'ha9; 
ram[16'h1110] = 8'hff; ram[16'h1111] = 8'h48; ram[16'h1112] = 8'ha9; ram[16'h1113] = 8'h37; ram[16'h1114] = 8'h28; ram[16'h1115] = 8'h73; ram[16'h1116] = 8'hea; ram[16'h1117] = 8'hea; 
ram[16'h1118] = 8'h08; ram[16'h1119] = 8'hc9; ram[16'h111a] = 8'h37; ram[16'h111b] = 8'hd0; ram[16'h111c] = 8'hfe; ram[16'h111d] = 8'h68; ram[16'h111e] = 8'h48; ram[16'h111f] = 8'hc9; 

ram[16'h1120] = 8'hff; ram[16'h1121] = 8'hd0; ram[16'h1122] = 8'hfe; ram[16'h1123] = 8'h28; ram[16'h1124] = 8'hc0; ram[16'h1125] = 8'h42; ram[16'h1126] = 8'hd0; ram[16'h1127] = 8'hfe; 
ram[16'h1128] = 8'he0; ram[16'h1129] = 8'h00; ram[16'h112a] = 8'hd0; ram[16'h112b] = 8'hfe; ram[16'h112c] = 8'ha0; ram[16'h112d] = 8'h42; ram[16'h112e] = 8'ha2; ram[16'h112f] = 8'h03; 
ram[16'h1130] = 8'h83; ram[16'h1131] = 8'hca; ram[16'h1132] = 8'hca; ram[16'h1133] = 8'hca; ram[16'h1134] = 8'hd0; ram[16'h1135] = 8'hfe; ram[16'h1136] = 8'ha9; ram[16'h1137] = 8'h00; 
ram[16'h1138] = 8'h48; ram[16'h1139] = 8'ha9; ram[16'h113a] = 8'h7c; ram[16'h113b] = 8'h28; ram[16'h113c] = 8'h83; ram[16'h113d] = 8'hea; ram[16'h113e] = 8'hea; ram[16'h113f] = 8'h08; 

ram[16'h1140] = 8'hc9; ram[16'h1141] = 8'h7c; ram[16'h1142] = 8'hd0; ram[16'h1143] = 8'hfe; ram[16'h1144] = 8'h68; ram[16'h1145] = 8'h48; ram[16'h1146] = 8'hc9; ram[16'h1147] = 8'h30; 
ram[16'h1148] = 8'hd0; ram[16'h1149] = 8'hfe; ram[16'h114a] = 8'h28; ram[16'h114b] = 8'ha9; ram[16'h114c] = 8'hff; ram[16'h114d] = 8'h48; ram[16'h114e] = 8'ha9; ram[16'h114f] = 8'h27; 
ram[16'h1150] = 8'h28; ram[16'h1151] = 8'h83; ram[16'h1152] = 8'hea; ram[16'h1153] = 8'hea; ram[16'h1154] = 8'h08; ram[16'h1155] = 8'hc9; ram[16'h1156] = 8'h27; ram[16'h1157] = 8'hd0; 
ram[16'h1158] = 8'hfe; ram[16'h1159] = 8'h68; ram[16'h115a] = 8'h48; ram[16'h115b] = 8'hc9; ram[16'h115c] = 8'hff; ram[16'h115d] = 8'hd0; ram[16'h115e] = 8'hfe; ram[16'h115f] = 8'h28; 

ram[16'h1160] = 8'hc0; ram[16'h1161] = 8'h42; ram[16'h1162] = 8'hd0; ram[16'h1163] = 8'hfe; ram[16'h1164] = 8'he0; ram[16'h1165] = 8'h00; ram[16'h1166] = 8'hd0; ram[16'h1167] = 8'hfe; 
ram[16'h1168] = 8'ha0; ram[16'h1169] = 8'h42; ram[16'h116a] = 8'ha2; ram[16'h116b] = 8'h03; ram[16'h116c] = 8'h93; ram[16'h116d] = 8'hca; ram[16'h116e] = 8'hca; ram[16'h116f] = 8'hca; 
ram[16'h1170] = 8'hd0; ram[16'h1171] = 8'hfe; ram[16'h1172] = 8'ha9; ram[16'h1173] = 8'h00; ram[16'h1174] = 8'h48; ram[16'h1175] = 8'ha9; ram[16'h1176] = 8'h6c; ram[16'h1177] = 8'h28; 
ram[16'h1178] = 8'h93; ram[16'h1179] = 8'hea; ram[16'h117a] = 8'hea; ram[16'h117b] = 8'h08; ram[16'h117c] = 8'hc9; ram[16'h117d] = 8'h6c; ram[16'h117e] = 8'hd0; ram[16'h117f] = 8'hfe; 

ram[16'h1180] = 8'h68; ram[16'h1181] = 8'h48; ram[16'h1182] = 8'hc9; ram[16'h1183] = 8'h30; ram[16'h1184] = 8'hd0; ram[16'h1185] = 8'hfe; ram[16'h1186] = 8'h28; ram[16'h1187] = 8'ha9; 
ram[16'h1188] = 8'hff; ram[16'h1189] = 8'h48; ram[16'h118a] = 8'ha9; ram[16'h118b] = 8'h17; ram[16'h118c] = 8'h28; ram[16'h118d] = 8'h93; ram[16'h118e] = 8'hea; ram[16'h118f] = 8'hea; 
ram[16'h1190] = 8'h08; ram[16'h1191] = 8'hc9; ram[16'h1192] = 8'h17; ram[16'h1193] = 8'hd0; ram[16'h1194] = 8'hfe; ram[16'h1195] = 8'h68; ram[16'h1196] = 8'h48; ram[16'h1197] = 8'hc9; 
ram[16'h1198] = 8'hff; ram[16'h1199] = 8'hd0; ram[16'h119a] = 8'hfe; ram[16'h119b] = 8'h28; ram[16'h119c] = 8'hc0; ram[16'h119d] = 8'h42; ram[16'h119e] = 8'hd0; ram[16'h119f] = 8'hfe; 

ram[16'h11a0] = 8'he0; ram[16'h11a1] = 8'h00; ram[16'h11a2] = 8'hd0; ram[16'h11a3] = 8'hfe; ram[16'h11a4] = 8'ha0; ram[16'h11a5] = 8'h42; ram[16'h11a6] = 8'ha2; ram[16'h11a7] = 8'h03; 
ram[16'h11a8] = 8'ha3; ram[16'h11a9] = 8'hca; ram[16'h11aa] = 8'hca; ram[16'h11ab] = 8'hca; ram[16'h11ac] = 8'hd0; ram[16'h11ad] = 8'hfe; ram[16'h11ae] = 8'ha9; ram[16'h11af] = 8'h00; 
ram[16'h11b0] = 8'h48; ram[16'h11b1] = 8'ha9; ram[16'h11b2] = 8'h5c; ram[16'h11b3] = 8'h28; ram[16'h11b4] = 8'ha3; ram[16'h11b5] = 8'hea; ram[16'h11b6] = 8'hea; ram[16'h11b7] = 8'h08; 
ram[16'h11b8] = 8'hc9; ram[16'h11b9] = 8'h5c; ram[16'h11ba] = 8'hd0; ram[16'h11bb] = 8'hfe; ram[16'h11bc] = 8'h68; ram[16'h11bd] = 8'h48; ram[16'h11be] = 8'hc9; ram[16'h11bf] = 8'h30; 

ram[16'h11c0] = 8'hd0; ram[16'h11c1] = 8'hfe; ram[16'h11c2] = 8'h28; ram[16'h11c3] = 8'ha9; ram[16'h11c4] = 8'hff; ram[16'h11c5] = 8'h48; ram[16'h11c6] = 8'ha9; ram[16'h11c7] = 8'h07; 
ram[16'h11c8] = 8'h28; ram[16'h11c9] = 8'ha3; ram[16'h11ca] = 8'hea; ram[16'h11cb] = 8'hea; ram[16'h11cc] = 8'h08; ram[16'h11cd] = 8'hc9; ram[16'h11ce] = 8'h07; ram[16'h11cf] = 8'hd0; 
ram[16'h11d0] = 8'hfe; ram[16'h11d1] = 8'h68; ram[16'h11d2] = 8'h48; ram[16'h11d3] = 8'hc9; ram[16'h11d4] = 8'hff; ram[16'h11d5] = 8'hd0; ram[16'h11d6] = 8'hfe; ram[16'h11d7] = 8'h28; 
ram[16'h11d8] = 8'hc0; ram[16'h11d9] = 8'h42; ram[16'h11da] = 8'hd0; ram[16'h11db] = 8'hfe; ram[16'h11dc] = 8'he0; ram[16'h11dd] = 8'h00; ram[16'h11de] = 8'hd0; ram[16'h11df] = 8'hfe; 

ram[16'h11e0] = 8'ha0; ram[16'h11e1] = 8'h42; ram[16'h11e2] = 8'ha2; ram[16'h11e3] = 8'h03; ram[16'h11e4] = 8'hb3; ram[16'h11e5] = 8'hca; ram[16'h11e6] = 8'hca; ram[16'h11e7] = 8'hca; 
ram[16'h11e8] = 8'hd0; ram[16'h11e9] = 8'hfe; ram[16'h11ea] = 8'ha9; ram[16'h11eb] = 8'h00; ram[16'h11ec] = 8'h48; ram[16'h11ed] = 8'ha9; ram[16'h11ee] = 8'h4c; ram[16'h11ef] = 8'h28; 
ram[16'h11f0] = 8'hb3; ram[16'h11f1] = 8'hea; ram[16'h11f2] = 8'hea; ram[16'h11f3] = 8'h08; ram[16'h11f4] = 8'hc9; ram[16'h11f5] = 8'h4c; ram[16'h11f6] = 8'hd0; ram[16'h11f7] = 8'hfe; 
ram[16'h11f8] = 8'h68; ram[16'h11f9] = 8'h48; ram[16'h11fa] = 8'hc9; ram[16'h11fb] = 8'h30; ram[16'h11fc] = 8'hd0; ram[16'h11fd] = 8'hfe; ram[16'h11fe] = 8'h28; ram[16'h11ff] = 8'ha9; 

ram[16'h1200] = 8'hff; ram[16'h1201] = 8'h48; ram[16'h1202] = 8'ha9; ram[16'h1203] = 8'hf7; ram[16'h1204] = 8'h28; ram[16'h1205] = 8'hb3; ram[16'h1206] = 8'hea; ram[16'h1207] = 8'hea; 
ram[16'h1208] = 8'h08; ram[16'h1209] = 8'hc9; ram[16'h120a] = 8'hf7; ram[16'h120b] = 8'hd0; ram[16'h120c] = 8'hfe; ram[16'h120d] = 8'h68; ram[16'h120e] = 8'h48; ram[16'h120f] = 8'hc9; 
ram[16'h1210] = 8'hff; ram[16'h1211] = 8'hd0; ram[16'h1212] = 8'hfe; ram[16'h1213] = 8'h28; ram[16'h1214] = 8'hc0; ram[16'h1215] = 8'h42; ram[16'h1216] = 8'hd0; ram[16'h1217] = 8'hfe; 
ram[16'h1218] = 8'he0; ram[16'h1219] = 8'h00; ram[16'h121a] = 8'hd0; ram[16'h121b] = 8'hfe; ram[16'h121c] = 8'ha0; ram[16'h121d] = 8'h42; ram[16'h121e] = 8'ha2; ram[16'h121f] = 8'h03; 

ram[16'h1220] = 8'hc3; ram[16'h1221] = 8'hca; ram[16'h1222] = 8'hca; ram[16'h1223] = 8'hca; ram[16'h1224] = 8'hd0; ram[16'h1225] = 8'hfe; ram[16'h1226] = 8'ha9; ram[16'h1227] = 8'h00; 
ram[16'h1228] = 8'h48; ram[16'h1229] = 8'ha9; ram[16'h122a] = 8'h3c; ram[16'h122b] = 8'h28; ram[16'h122c] = 8'hc3; ram[16'h122d] = 8'hea; ram[16'h122e] = 8'hea; ram[16'h122f] = 8'h08; 
ram[16'h1230] = 8'hc9; ram[16'h1231] = 8'h3c; ram[16'h1232] = 8'hd0; ram[16'h1233] = 8'hfe; ram[16'h1234] = 8'h68; ram[16'h1235] = 8'h48; ram[16'h1236] = 8'hc9; ram[16'h1237] = 8'h30; 
ram[16'h1238] = 8'hd0; ram[16'h1239] = 8'hfe; ram[16'h123a] = 8'h28; ram[16'h123b] = 8'ha9; ram[16'h123c] = 8'hff; ram[16'h123d] = 8'h48; ram[16'h123e] = 8'ha9; ram[16'h123f] = 8'he7; 

ram[16'h1240] = 8'h28; ram[16'h1241] = 8'hc3; ram[16'h1242] = 8'hea; ram[16'h1243] = 8'hea; ram[16'h1244] = 8'h08; ram[16'h1245] = 8'hc9; ram[16'h1246] = 8'he7; ram[16'h1247] = 8'hd0; 
ram[16'h1248] = 8'hfe; ram[16'h1249] = 8'h68; ram[16'h124a] = 8'h48; ram[16'h124b] = 8'hc9; ram[16'h124c] = 8'hff; ram[16'h124d] = 8'hd0; ram[16'h124e] = 8'hfe; ram[16'h124f] = 8'h28; 
ram[16'h1250] = 8'hc0; ram[16'h1251] = 8'h42; ram[16'h1252] = 8'hd0; ram[16'h1253] = 8'hfe; ram[16'h1254] = 8'he0; ram[16'h1255] = 8'h00; ram[16'h1256] = 8'hd0; ram[16'h1257] = 8'hfe; 
ram[16'h1258] = 8'ha0; ram[16'h1259] = 8'h42; ram[16'h125a] = 8'ha2; ram[16'h125b] = 8'h03; ram[16'h125c] = 8'hd3; ram[16'h125d] = 8'hca; ram[16'h125e] = 8'hca; ram[16'h125f] = 8'hca; 

ram[16'h1260] = 8'hd0; ram[16'h1261] = 8'hfe; ram[16'h1262] = 8'ha9; ram[16'h1263] = 8'h00; ram[16'h1264] = 8'h48; ram[16'h1265] = 8'ha9; ram[16'h1266] = 8'h2c; ram[16'h1267] = 8'h28; 
ram[16'h1268] = 8'hd3; ram[16'h1269] = 8'hea; ram[16'h126a] = 8'hea; ram[16'h126b] = 8'h08; ram[16'h126c] = 8'hc9; ram[16'h126d] = 8'h2c; ram[16'h126e] = 8'hd0; ram[16'h126f] = 8'hfe; 
ram[16'h1270] = 8'h68; ram[16'h1271] = 8'h48; ram[16'h1272] = 8'hc9; ram[16'h1273] = 8'h30; ram[16'h1274] = 8'hd0; ram[16'h1275] = 8'hfe; ram[16'h1276] = 8'h28; ram[16'h1277] = 8'ha9; 
ram[16'h1278] = 8'hff; ram[16'h1279] = 8'h48; ram[16'h127a] = 8'ha9; ram[16'h127b] = 8'hd7; ram[16'h127c] = 8'h28; ram[16'h127d] = 8'hd3; ram[16'h127e] = 8'hea; ram[16'h127f] = 8'hea; 

ram[16'h1280] = 8'h08; ram[16'h1281] = 8'hc9; ram[16'h1282] = 8'hd7; ram[16'h1283] = 8'hd0; ram[16'h1284] = 8'hfe; ram[16'h1285] = 8'h68; ram[16'h1286] = 8'h48; ram[16'h1287] = 8'hc9; 
ram[16'h1288] = 8'hff; ram[16'h1289] = 8'hd0; ram[16'h128a] = 8'hfe; ram[16'h128b] = 8'h28; ram[16'h128c] = 8'hc0; ram[16'h128d] = 8'h42; ram[16'h128e] = 8'hd0; ram[16'h128f] = 8'hfe; 
ram[16'h1290] = 8'he0; ram[16'h1291] = 8'h00; ram[16'h1292] = 8'hd0; ram[16'h1293] = 8'hfe; ram[16'h1294] = 8'ha0; ram[16'h1295] = 8'h42; ram[16'h1296] = 8'ha2; ram[16'h1297] = 8'h03; 
ram[16'h1298] = 8'he3; ram[16'h1299] = 8'hca; ram[16'h129a] = 8'hca; ram[16'h129b] = 8'hca; ram[16'h129c] = 8'hd0; ram[16'h129d] = 8'hfe; ram[16'h129e] = 8'ha9; ram[16'h129f] = 8'h00; 

ram[16'h12a0] = 8'h48; ram[16'h12a1] = 8'ha9; ram[16'h12a2] = 8'h1c; ram[16'h12a3] = 8'h28; ram[16'h12a4] = 8'he3; ram[16'h12a5] = 8'hea; ram[16'h12a6] = 8'hea; ram[16'h12a7] = 8'h08; 
ram[16'h12a8] = 8'hc9; ram[16'h12a9] = 8'h1c; ram[16'h12aa] = 8'hd0; ram[16'h12ab] = 8'hfe; ram[16'h12ac] = 8'h68; ram[16'h12ad] = 8'h48; ram[16'h12ae] = 8'hc9; ram[16'h12af] = 8'h30; 
ram[16'h12b0] = 8'hd0; ram[16'h12b1] = 8'hfe; ram[16'h12b2] = 8'h28; ram[16'h12b3] = 8'ha9; ram[16'h12b4] = 8'hff; ram[16'h12b5] = 8'h48; ram[16'h12b6] = 8'ha9; ram[16'h12b7] = 8'hc7; 
ram[16'h12b8] = 8'h28; ram[16'h12b9] = 8'he3; ram[16'h12ba] = 8'hea; ram[16'h12bb] = 8'hea; ram[16'h12bc] = 8'h08; ram[16'h12bd] = 8'hc9; ram[16'h12be] = 8'hc7; ram[16'h12bf] = 8'hd0; 

ram[16'h12c0] = 8'hfe; ram[16'h12c1] = 8'h68; ram[16'h12c2] = 8'h48; ram[16'h12c3] = 8'hc9; ram[16'h12c4] = 8'hff; ram[16'h12c5] = 8'hd0; ram[16'h12c6] = 8'hfe; ram[16'h12c7] = 8'h28; 
ram[16'h12c8] = 8'hc0; ram[16'h12c9] = 8'h42; ram[16'h12ca] = 8'hd0; ram[16'h12cb] = 8'hfe; ram[16'h12cc] = 8'he0; ram[16'h12cd] = 8'h00; ram[16'h12ce] = 8'hd0; ram[16'h12cf] = 8'hfe; 
ram[16'h12d0] = 8'ha0; ram[16'h12d1] = 8'h42; ram[16'h12d2] = 8'ha2; ram[16'h12d3] = 8'h03; ram[16'h12d4] = 8'hf3; ram[16'h12d5] = 8'hca; ram[16'h12d6] = 8'hca; ram[16'h12d7] = 8'hca; 
ram[16'h12d8] = 8'hd0; ram[16'h12d9] = 8'hfe; ram[16'h12da] = 8'ha9; ram[16'h12db] = 8'h00; ram[16'h12dc] = 8'h48; ram[16'h12dd] = 8'ha9; ram[16'h12de] = 8'h0c; ram[16'h12df] = 8'h28; 

ram[16'h12e0] = 8'hf3; ram[16'h12e1] = 8'hea; ram[16'h12e2] = 8'hea; ram[16'h12e3] = 8'h08; ram[16'h12e4] = 8'hc9; ram[16'h12e5] = 8'h0c; ram[16'h12e6] = 8'hd0; ram[16'h12e7] = 8'hfe; 
ram[16'h12e8] = 8'h68; ram[16'h12e9] = 8'h48; ram[16'h12ea] = 8'hc9; ram[16'h12eb] = 8'h30; ram[16'h12ec] = 8'hd0; ram[16'h12ed] = 8'hfe; ram[16'h12ee] = 8'h28; ram[16'h12ef] = 8'ha9; 
ram[16'h12f0] = 8'hff; ram[16'h12f1] = 8'h48; ram[16'h12f2] = 8'ha9; ram[16'h12f3] = 8'hb7; ram[16'h12f4] = 8'h28; ram[16'h12f5] = 8'hf3; ram[16'h12f6] = 8'hea; ram[16'h12f7] = 8'hea; 
ram[16'h12f8] = 8'h08; ram[16'h12f9] = 8'hc9; ram[16'h12fa] = 8'hb7; ram[16'h12fb] = 8'hd0; ram[16'h12fc] = 8'hfe; ram[16'h12fd] = 8'h68; ram[16'h12fe] = 8'h48; ram[16'h12ff] = 8'hc9; 

ram[16'h1300] = 8'hff; ram[16'h1301] = 8'hd0; ram[16'h1302] = 8'hfe; ram[16'h1303] = 8'h28; ram[16'h1304] = 8'hc0; ram[16'h1305] = 8'h42; ram[16'h1306] = 8'hd0; ram[16'h1307] = 8'hfe; 
ram[16'h1308] = 8'he0; ram[16'h1309] = 8'h00; ram[16'h130a] = 8'hd0; ram[16'h130b] = 8'hfe; ram[16'h130c] = 8'ha0; ram[16'h130d] = 8'h42; ram[16'h130e] = 8'ha2; ram[16'h130f] = 8'h03; 
ram[16'h1310] = 8'h0b; ram[16'h1311] = 8'hca; ram[16'h1312] = 8'hca; ram[16'h1313] = 8'hca; ram[16'h1314] = 8'hd0; ram[16'h1315] = 8'hfe; ram[16'h1316] = 8'ha9; ram[16'h1317] = 8'h00; 
ram[16'h1318] = 8'h48; ram[16'h1319] = 8'ha9; ram[16'h131a] = 8'hf4; ram[16'h131b] = 8'h28; ram[16'h131c] = 8'h0b; ram[16'h131d] = 8'hea; ram[16'h131e] = 8'hea; ram[16'h131f] = 8'h08; 

ram[16'h1320] = 8'hc9; ram[16'h1321] = 8'hf4; ram[16'h1322] = 8'hd0; ram[16'h1323] = 8'hfe; ram[16'h1324] = 8'h68; ram[16'h1325] = 8'h48; ram[16'h1326] = 8'hc9; ram[16'h1327] = 8'h30; 
ram[16'h1328] = 8'hd0; ram[16'h1329] = 8'hfe; ram[16'h132a] = 8'h28; ram[16'h132b] = 8'ha9; ram[16'h132c] = 8'hff; ram[16'h132d] = 8'h48; ram[16'h132e] = 8'ha9; ram[16'h132f] = 8'h9f; 
ram[16'h1330] = 8'h28; ram[16'h1331] = 8'h0b; ram[16'h1332] = 8'hea; ram[16'h1333] = 8'hea; ram[16'h1334] = 8'h08; ram[16'h1335] = 8'hc9; ram[16'h1336] = 8'h9f; ram[16'h1337] = 8'hd0; 
ram[16'h1338] = 8'hfe; ram[16'h1339] = 8'h68; ram[16'h133a] = 8'h48; ram[16'h133b] = 8'hc9; ram[16'h133c] = 8'hff; ram[16'h133d] = 8'hd0; ram[16'h133e] = 8'hfe; ram[16'h133f] = 8'h28; 

ram[16'h1340] = 8'hc0; ram[16'h1341] = 8'h42; ram[16'h1342] = 8'hd0; ram[16'h1343] = 8'hfe; ram[16'h1344] = 8'he0; ram[16'h1345] = 8'h00; ram[16'h1346] = 8'hd0; ram[16'h1347] = 8'hfe; 
ram[16'h1348] = 8'ha0; ram[16'h1349] = 8'h42; ram[16'h134a] = 8'ha2; ram[16'h134b] = 8'h03; ram[16'h134c] = 8'h1b; ram[16'h134d] = 8'hca; ram[16'h134e] = 8'hca; ram[16'h134f] = 8'hca; 
ram[16'h1350] = 8'hd0; ram[16'h1351] = 8'hfe; ram[16'h1352] = 8'ha9; ram[16'h1353] = 8'h00; ram[16'h1354] = 8'h48; ram[16'h1355] = 8'ha9; ram[16'h1356] = 8'he4; ram[16'h1357] = 8'h28; 
ram[16'h1358] = 8'h1b; ram[16'h1359] = 8'hea; ram[16'h135a] = 8'hea; ram[16'h135b] = 8'h08; ram[16'h135c] = 8'hc9; ram[16'h135d] = 8'he4; ram[16'h135e] = 8'hd0; ram[16'h135f] = 8'hfe; 

ram[16'h1360] = 8'h68; ram[16'h1361] = 8'h48; ram[16'h1362] = 8'hc9; ram[16'h1363] = 8'h30; ram[16'h1364] = 8'hd0; ram[16'h1365] = 8'hfe; ram[16'h1366] = 8'h28; ram[16'h1367] = 8'ha9; 
ram[16'h1368] = 8'hff; ram[16'h1369] = 8'h48; ram[16'h136a] = 8'ha9; ram[16'h136b] = 8'h8f; ram[16'h136c] = 8'h28; ram[16'h136d] = 8'h1b; ram[16'h136e] = 8'hea; ram[16'h136f] = 8'hea; 
ram[16'h1370] = 8'h08; ram[16'h1371] = 8'hc9; ram[16'h1372] = 8'h8f; ram[16'h1373] = 8'hd0; ram[16'h1374] = 8'hfe; ram[16'h1375] = 8'h68; ram[16'h1376] = 8'h48; ram[16'h1377] = 8'hc9; 
ram[16'h1378] = 8'hff; ram[16'h1379] = 8'hd0; ram[16'h137a] = 8'hfe; ram[16'h137b] = 8'h28; ram[16'h137c] = 8'hc0; ram[16'h137d] = 8'h42; ram[16'h137e] = 8'hd0; ram[16'h137f] = 8'hfe; 

ram[16'h1380] = 8'he0; ram[16'h1381] = 8'h00; ram[16'h1382] = 8'hd0; ram[16'h1383] = 8'hfe; ram[16'h1384] = 8'ha0; ram[16'h1385] = 8'h42; ram[16'h1386] = 8'ha2; ram[16'h1387] = 8'h03; 
ram[16'h1388] = 8'h2b; ram[16'h1389] = 8'hca; ram[16'h138a] = 8'hca; ram[16'h138b] = 8'hca; ram[16'h138c] = 8'hd0; ram[16'h138d] = 8'hfe; ram[16'h138e] = 8'ha9; ram[16'h138f] = 8'h00; 
ram[16'h1390] = 8'h48; ram[16'h1391] = 8'ha9; ram[16'h1392] = 8'hd4; ram[16'h1393] = 8'h28; ram[16'h1394] = 8'h2b; ram[16'h1395] = 8'hea; ram[16'h1396] = 8'hea; ram[16'h1397] = 8'h08; 
ram[16'h1398] = 8'hc9; ram[16'h1399] = 8'hd4; ram[16'h139a] = 8'hd0; ram[16'h139b] = 8'hfe; ram[16'h139c] = 8'h68; ram[16'h139d] = 8'h48; ram[16'h139e] = 8'hc9; ram[16'h139f] = 8'h30; 

ram[16'h13a0] = 8'hd0; ram[16'h13a1] = 8'hfe; ram[16'h13a2] = 8'h28; ram[16'h13a3] = 8'ha9; ram[16'h13a4] = 8'hff; ram[16'h13a5] = 8'h48; ram[16'h13a6] = 8'ha9; ram[16'h13a7] = 8'h7f; 
ram[16'h13a8] = 8'h28; ram[16'h13a9] = 8'h2b; ram[16'h13aa] = 8'hea; ram[16'h13ab] = 8'hea; ram[16'h13ac] = 8'h08; ram[16'h13ad] = 8'hc9; ram[16'h13ae] = 8'h7f; ram[16'h13af] = 8'hd0; 
ram[16'h13b0] = 8'hfe; ram[16'h13b1] = 8'h68; ram[16'h13b2] = 8'h48; ram[16'h13b3] = 8'hc9; ram[16'h13b4] = 8'hff; ram[16'h13b5] = 8'hd0; ram[16'h13b6] = 8'hfe; ram[16'h13b7] = 8'h28; 
ram[16'h13b8] = 8'hc0; ram[16'h13b9] = 8'h42; ram[16'h13ba] = 8'hd0; ram[16'h13bb] = 8'hfe; ram[16'h13bc] = 8'he0; ram[16'h13bd] = 8'h00; ram[16'h13be] = 8'hd0; ram[16'h13bf] = 8'hfe; 

ram[16'h13c0] = 8'ha0; ram[16'h13c1] = 8'h42; ram[16'h13c2] = 8'ha2; ram[16'h13c3] = 8'h03; ram[16'h13c4] = 8'h3b; ram[16'h13c5] = 8'hca; ram[16'h13c6] = 8'hca; ram[16'h13c7] = 8'hca; 
ram[16'h13c8] = 8'hd0; ram[16'h13c9] = 8'hfe; ram[16'h13ca] = 8'ha9; ram[16'h13cb] = 8'h00; ram[16'h13cc] = 8'h48; ram[16'h13cd] = 8'ha9; ram[16'h13ce] = 8'hc4; ram[16'h13cf] = 8'h28; 
ram[16'h13d0] = 8'h3b; ram[16'h13d1] = 8'hea; ram[16'h13d2] = 8'hea; ram[16'h13d3] = 8'h08; ram[16'h13d4] = 8'hc9; ram[16'h13d5] = 8'hc4; ram[16'h13d6] = 8'hd0; ram[16'h13d7] = 8'hfe; 
ram[16'h13d8] = 8'h68; ram[16'h13d9] = 8'h48; ram[16'h13da] = 8'hc9; ram[16'h13db] = 8'h30; ram[16'h13dc] = 8'hd0; ram[16'h13dd] = 8'hfe; ram[16'h13de] = 8'h28; ram[16'h13df] = 8'ha9; 

ram[16'h13e0] = 8'hff; ram[16'h13e1] = 8'h48; ram[16'h13e2] = 8'ha9; ram[16'h13e3] = 8'h6f; ram[16'h13e4] = 8'h28; ram[16'h13e5] = 8'h3b; ram[16'h13e6] = 8'hea; ram[16'h13e7] = 8'hea; 
ram[16'h13e8] = 8'h08; ram[16'h13e9] = 8'hc9; ram[16'h13ea] = 8'h6f; ram[16'h13eb] = 8'hd0; ram[16'h13ec] = 8'hfe; ram[16'h13ed] = 8'h68; ram[16'h13ee] = 8'h48; ram[16'h13ef] = 8'hc9; 
ram[16'h13f0] = 8'hff; ram[16'h13f1] = 8'hd0; ram[16'h13f2] = 8'hfe; ram[16'h13f3] = 8'h28; ram[16'h13f4] = 8'hc0; ram[16'h13f5] = 8'h42; ram[16'h13f6] = 8'hd0; ram[16'h13f7] = 8'hfe; 
ram[16'h13f8] = 8'he0; ram[16'h13f9] = 8'h00; ram[16'h13fa] = 8'hd0; ram[16'h13fb] = 8'hfe; ram[16'h13fc] = 8'ha0; ram[16'h13fd] = 8'h42; ram[16'h13fe] = 8'ha2; ram[16'h13ff] = 8'h03; 

ram[16'h1400] = 8'h4b; ram[16'h1401] = 8'hca; ram[16'h1402] = 8'hca; ram[16'h1403] = 8'hca; ram[16'h1404] = 8'hd0; ram[16'h1405] = 8'hfe; ram[16'h1406] = 8'ha9; ram[16'h1407] = 8'h00; 
ram[16'h1408] = 8'h48; ram[16'h1409] = 8'ha9; ram[16'h140a] = 8'hb4; ram[16'h140b] = 8'h28; ram[16'h140c] = 8'h4b; ram[16'h140d] = 8'hea; ram[16'h140e] = 8'hea; ram[16'h140f] = 8'h08; 
ram[16'h1410] = 8'hc9; ram[16'h1411] = 8'hb4; ram[16'h1412] = 8'hd0; ram[16'h1413] = 8'hfe; ram[16'h1414] = 8'h68; ram[16'h1415] = 8'h48; ram[16'h1416] = 8'hc9; ram[16'h1417] = 8'h30; 
ram[16'h1418] = 8'hd0; ram[16'h1419] = 8'hfe; ram[16'h141a] = 8'h28; ram[16'h141b] = 8'ha9; ram[16'h141c] = 8'hff; ram[16'h141d] = 8'h48; ram[16'h141e] = 8'ha9; ram[16'h141f] = 8'h5f; 

ram[16'h1420] = 8'h28; ram[16'h1421] = 8'h4b; ram[16'h1422] = 8'hea; ram[16'h1423] = 8'hea; ram[16'h1424] = 8'h08; ram[16'h1425] = 8'hc9; ram[16'h1426] = 8'h5f; ram[16'h1427] = 8'hd0; 
ram[16'h1428] = 8'hfe; ram[16'h1429] = 8'h68; ram[16'h142a] = 8'h48; ram[16'h142b] = 8'hc9; ram[16'h142c] = 8'hff; ram[16'h142d] = 8'hd0; ram[16'h142e] = 8'hfe; ram[16'h142f] = 8'h28; 
ram[16'h1430] = 8'hc0; ram[16'h1431] = 8'h42; ram[16'h1432] = 8'hd0; ram[16'h1433] = 8'hfe; ram[16'h1434] = 8'he0; ram[16'h1435] = 8'h00; ram[16'h1436] = 8'hd0; ram[16'h1437] = 8'hfe; 
ram[16'h1438] = 8'ha0; ram[16'h1439] = 8'h42; ram[16'h143a] = 8'ha2; ram[16'h143b] = 8'h03; ram[16'h143c] = 8'h5b; ram[16'h143d] = 8'hca; ram[16'h143e] = 8'hca; ram[16'h143f] = 8'hca; 

ram[16'h1440] = 8'hd0; ram[16'h1441] = 8'hfe; ram[16'h1442] = 8'ha9; ram[16'h1443] = 8'h00; ram[16'h1444] = 8'h48; ram[16'h1445] = 8'ha9; ram[16'h1446] = 8'ha4; ram[16'h1447] = 8'h28; 
ram[16'h1448] = 8'h5b; ram[16'h1449] = 8'hea; ram[16'h144a] = 8'hea; ram[16'h144b] = 8'h08; ram[16'h144c] = 8'hc9; ram[16'h144d] = 8'ha4; ram[16'h144e] = 8'hd0; ram[16'h144f] = 8'hfe; 
ram[16'h1450] = 8'h68; ram[16'h1451] = 8'h48; ram[16'h1452] = 8'hc9; ram[16'h1453] = 8'h30; ram[16'h1454] = 8'hd0; ram[16'h1455] = 8'hfe; ram[16'h1456] = 8'h28; ram[16'h1457] = 8'ha9; 
ram[16'h1458] = 8'hff; ram[16'h1459] = 8'h48; ram[16'h145a] = 8'ha9; ram[16'h145b] = 8'h4f; ram[16'h145c] = 8'h28; ram[16'h145d] = 8'h5b; ram[16'h145e] = 8'hea; ram[16'h145f] = 8'hea; 

ram[16'h1460] = 8'h08; ram[16'h1461] = 8'hc9; ram[16'h1462] = 8'h4f; ram[16'h1463] = 8'hd0; ram[16'h1464] = 8'hfe; ram[16'h1465] = 8'h68; ram[16'h1466] = 8'h48; ram[16'h1467] = 8'hc9; 
ram[16'h1468] = 8'hff; ram[16'h1469] = 8'hd0; ram[16'h146a] = 8'hfe; ram[16'h146b] = 8'h28; ram[16'h146c] = 8'hc0; ram[16'h146d] = 8'h42; ram[16'h146e] = 8'hd0; ram[16'h146f] = 8'hfe; 
ram[16'h1470] = 8'he0; ram[16'h1471] = 8'h00; ram[16'h1472] = 8'hd0; ram[16'h1473] = 8'hfe; ram[16'h1474] = 8'ha0; ram[16'h1475] = 8'h42; ram[16'h1476] = 8'ha2; ram[16'h1477] = 8'h03; 
ram[16'h1478] = 8'h6b; ram[16'h1479] = 8'hca; ram[16'h147a] = 8'hca; ram[16'h147b] = 8'hca; ram[16'h147c] = 8'hd0; ram[16'h147d] = 8'hfe; ram[16'h147e] = 8'ha9; ram[16'h147f] = 8'h00; 

ram[16'h1480] = 8'h48; ram[16'h1481] = 8'ha9; ram[16'h1482] = 8'h94; ram[16'h1483] = 8'h28; ram[16'h1484] = 8'h6b; ram[16'h1485] = 8'hea; ram[16'h1486] = 8'hea; ram[16'h1487] = 8'h08; 
ram[16'h1488] = 8'hc9; ram[16'h1489] = 8'h94; ram[16'h148a] = 8'hd0; ram[16'h148b] = 8'hfe; ram[16'h148c] = 8'h68; ram[16'h148d] = 8'h48; ram[16'h148e] = 8'hc9; ram[16'h148f] = 8'h30; 
ram[16'h1490] = 8'hd0; ram[16'h1491] = 8'hfe; ram[16'h1492] = 8'h28; ram[16'h1493] = 8'ha9; ram[16'h1494] = 8'hff; ram[16'h1495] = 8'h48; ram[16'h1496] = 8'ha9; ram[16'h1497] = 8'h3f; 
ram[16'h1498] = 8'h28; ram[16'h1499] = 8'h6b; ram[16'h149a] = 8'hea; ram[16'h149b] = 8'hea; ram[16'h149c] = 8'h08; ram[16'h149d] = 8'hc9; ram[16'h149e] = 8'h3f; ram[16'h149f] = 8'hd0; 

ram[16'h14a0] = 8'hfe; ram[16'h14a1] = 8'h68; ram[16'h14a2] = 8'h48; ram[16'h14a3] = 8'hc9; ram[16'h14a4] = 8'hff; ram[16'h14a5] = 8'hd0; ram[16'h14a6] = 8'hfe; ram[16'h14a7] = 8'h28; 
ram[16'h14a8] = 8'hc0; ram[16'h14a9] = 8'h42; ram[16'h14aa] = 8'hd0; ram[16'h14ab] = 8'hfe; ram[16'h14ac] = 8'he0; ram[16'h14ad] = 8'h00; ram[16'h14ae] = 8'hd0; ram[16'h14af] = 8'hfe; 
ram[16'h14b0] = 8'ha0; ram[16'h14b1] = 8'h42; ram[16'h14b2] = 8'ha2; ram[16'h14b3] = 8'h03; ram[16'h14b4] = 8'h7b; ram[16'h14b5] = 8'hca; ram[16'h14b6] = 8'hca; ram[16'h14b7] = 8'hca; 
ram[16'h14b8] = 8'hd0; ram[16'h14b9] = 8'hfe; ram[16'h14ba] = 8'ha9; ram[16'h14bb] = 8'h00; ram[16'h14bc] = 8'h48; ram[16'h14bd] = 8'ha9; ram[16'h14be] = 8'h84; ram[16'h14bf] = 8'h28; 

ram[16'h14c0] = 8'h7b; ram[16'h14c1] = 8'hea; ram[16'h14c2] = 8'hea; ram[16'h14c3] = 8'h08; ram[16'h14c4] = 8'hc9; ram[16'h14c5] = 8'h84; ram[16'h14c6] = 8'hd0; ram[16'h14c7] = 8'hfe; 
ram[16'h14c8] = 8'h68; ram[16'h14c9] = 8'h48; ram[16'h14ca] = 8'hc9; ram[16'h14cb] = 8'h30; ram[16'h14cc] = 8'hd0; ram[16'h14cd] = 8'hfe; ram[16'h14ce] = 8'h28; ram[16'h14cf] = 8'ha9; 
ram[16'h14d0] = 8'hff; ram[16'h14d1] = 8'h48; ram[16'h14d2] = 8'ha9; ram[16'h14d3] = 8'h2f; ram[16'h14d4] = 8'h28; ram[16'h14d5] = 8'h7b; ram[16'h14d6] = 8'hea; ram[16'h14d7] = 8'hea; 
ram[16'h14d8] = 8'h08; ram[16'h14d9] = 8'hc9; ram[16'h14da] = 8'h2f; ram[16'h14db] = 8'hd0; ram[16'h14dc] = 8'hfe; ram[16'h14dd] = 8'h68; ram[16'h14de] = 8'h48; ram[16'h14df] = 8'hc9; 

ram[16'h14e0] = 8'hff; ram[16'h14e1] = 8'hd0; ram[16'h14e2] = 8'hfe; ram[16'h14e3] = 8'h28; ram[16'h14e4] = 8'hc0; ram[16'h14e5] = 8'h42; ram[16'h14e6] = 8'hd0; ram[16'h14e7] = 8'hfe; 
ram[16'h14e8] = 8'he0; ram[16'h14e9] = 8'h00; ram[16'h14ea] = 8'hd0; ram[16'h14eb] = 8'hfe; ram[16'h14ec] = 8'ha0; ram[16'h14ed] = 8'h42; ram[16'h14ee] = 8'ha2; ram[16'h14ef] = 8'h03; 
ram[16'h14f0] = 8'h8b; ram[16'h14f1] = 8'hca; ram[16'h14f2] = 8'hca; ram[16'h14f3] = 8'hca; ram[16'h14f4] = 8'hd0; ram[16'h14f5] = 8'hfe; ram[16'h14f6] = 8'ha9; ram[16'h14f7] = 8'h00; 
ram[16'h14f8] = 8'h48; ram[16'h14f9] = 8'ha9; ram[16'h14fa] = 8'h74; ram[16'h14fb] = 8'h28; ram[16'h14fc] = 8'h8b; ram[16'h14fd] = 8'hea; ram[16'h14fe] = 8'hea; ram[16'h14ff] = 8'h08; 

ram[16'h1500] = 8'hc9; ram[16'h1501] = 8'h74; ram[16'h1502] = 8'hd0; ram[16'h1503] = 8'hfe; ram[16'h1504] = 8'h68; ram[16'h1505] = 8'h48; ram[16'h1506] = 8'hc9; ram[16'h1507] = 8'h30; 
ram[16'h1508] = 8'hd0; ram[16'h1509] = 8'hfe; ram[16'h150a] = 8'h28; ram[16'h150b] = 8'ha9; ram[16'h150c] = 8'hff; ram[16'h150d] = 8'h48; ram[16'h150e] = 8'ha9; ram[16'h150f] = 8'h1f; 
ram[16'h1510] = 8'h28; ram[16'h1511] = 8'h8b; ram[16'h1512] = 8'hea; ram[16'h1513] = 8'hea; ram[16'h1514] = 8'h08; ram[16'h1515] = 8'hc9; ram[16'h1516] = 8'h1f; ram[16'h1517] = 8'hd0; 
ram[16'h1518] = 8'hfe; ram[16'h1519] = 8'h68; ram[16'h151a] = 8'h48; ram[16'h151b] = 8'hc9; ram[16'h151c] = 8'hff; ram[16'h151d] = 8'hd0; ram[16'h151e] = 8'hfe; ram[16'h151f] = 8'h28; 

ram[16'h1520] = 8'hc0; ram[16'h1521] = 8'h42; ram[16'h1522] = 8'hd0; ram[16'h1523] = 8'hfe; ram[16'h1524] = 8'he0; ram[16'h1525] = 8'h00; ram[16'h1526] = 8'hd0; ram[16'h1527] = 8'hfe; 
ram[16'h1528] = 8'ha0; ram[16'h1529] = 8'h42; ram[16'h152a] = 8'ha2; ram[16'h152b] = 8'h03; ram[16'h152c] = 8'h9b; ram[16'h152d] = 8'hca; ram[16'h152e] = 8'hca; ram[16'h152f] = 8'hca; 
ram[16'h1530] = 8'hd0; ram[16'h1531] = 8'hfe; ram[16'h1532] = 8'ha9; ram[16'h1533] = 8'h00; ram[16'h1534] = 8'h48; ram[16'h1535] = 8'ha9; ram[16'h1536] = 8'h64; ram[16'h1537] = 8'h28; 
ram[16'h1538] = 8'h9b; ram[16'h1539] = 8'hea; ram[16'h153a] = 8'hea; ram[16'h153b] = 8'h08; ram[16'h153c] = 8'hc9; ram[16'h153d] = 8'h64; ram[16'h153e] = 8'hd0; ram[16'h153f] = 8'hfe; 

ram[16'h1540] = 8'h68; ram[16'h1541] = 8'h48; ram[16'h1542] = 8'hc9; ram[16'h1543] = 8'h30; ram[16'h1544] = 8'hd0; ram[16'h1545] = 8'hfe; ram[16'h1546] = 8'h28; ram[16'h1547] = 8'ha9; 
ram[16'h1548] = 8'hff; ram[16'h1549] = 8'h48; ram[16'h154a] = 8'ha9; ram[16'h154b] = 8'h0f; ram[16'h154c] = 8'h28; ram[16'h154d] = 8'h9b; ram[16'h154e] = 8'hea; ram[16'h154f] = 8'hea; 
ram[16'h1550] = 8'h08; ram[16'h1551] = 8'hc9; ram[16'h1552] = 8'h0f; ram[16'h1553] = 8'hd0; ram[16'h1554] = 8'hfe; ram[16'h1555] = 8'h68; ram[16'h1556] = 8'h48; ram[16'h1557] = 8'hc9; 
ram[16'h1558] = 8'hff; ram[16'h1559] = 8'hd0; ram[16'h155a] = 8'hfe; ram[16'h155b] = 8'h28; ram[16'h155c] = 8'hc0; ram[16'h155d] = 8'h42; ram[16'h155e] = 8'hd0; ram[16'h155f] = 8'hfe; 

ram[16'h1560] = 8'he0; ram[16'h1561] = 8'h00; ram[16'h1562] = 8'hd0; ram[16'h1563] = 8'hfe; ram[16'h1564] = 8'ha0; ram[16'h1565] = 8'h42; ram[16'h1566] = 8'ha2; ram[16'h1567] = 8'h03; 
ram[16'h1568] = 8'hab; ram[16'h1569] = 8'hca; ram[16'h156a] = 8'hca; ram[16'h156b] = 8'hca; ram[16'h156c] = 8'hd0; ram[16'h156d] = 8'hfe; ram[16'h156e] = 8'ha9; ram[16'h156f] = 8'h00; 
ram[16'h1570] = 8'h48; ram[16'h1571] = 8'ha9; ram[16'h1572] = 8'h54; ram[16'h1573] = 8'h28; ram[16'h1574] = 8'hab; ram[16'h1575] = 8'hea; ram[16'h1576] = 8'hea; ram[16'h1577] = 8'h08; 
ram[16'h1578] = 8'hc9; ram[16'h1579] = 8'h54; ram[16'h157a] = 8'hd0; ram[16'h157b] = 8'hfe; ram[16'h157c] = 8'h68; ram[16'h157d] = 8'h48; ram[16'h157e] = 8'hc9; ram[16'h157f] = 8'h30; 

ram[16'h1580] = 8'hd0; ram[16'h1581] = 8'hfe; ram[16'h1582] = 8'h28; ram[16'h1583] = 8'ha9; ram[16'h1584] = 8'hff; ram[16'h1585] = 8'h48; ram[16'h1586] = 8'ha9; ram[16'h1587] = 8'hff; 
ram[16'h1588] = 8'h28; ram[16'h1589] = 8'hab; ram[16'h158a] = 8'hea; ram[16'h158b] = 8'hea; ram[16'h158c] = 8'h08; ram[16'h158d] = 8'hc9; ram[16'h158e] = 8'hff; ram[16'h158f] = 8'hd0; 
ram[16'h1590] = 8'hfe; ram[16'h1591] = 8'h68; ram[16'h1592] = 8'h48; ram[16'h1593] = 8'hc9; ram[16'h1594] = 8'hff; ram[16'h1595] = 8'hd0; ram[16'h1596] = 8'hfe; ram[16'h1597] = 8'h28; 
ram[16'h1598] = 8'hc0; ram[16'h1599] = 8'h42; ram[16'h159a] = 8'hd0; ram[16'h159b] = 8'hfe; ram[16'h159c] = 8'he0; ram[16'h159d] = 8'h00; ram[16'h159e] = 8'hd0; ram[16'h159f] = 8'hfe; 

ram[16'h15a0] = 8'ha0; ram[16'h15a1] = 8'h42; ram[16'h15a2] = 8'ha2; ram[16'h15a3] = 8'h03; ram[16'h15a4] = 8'hbb; ram[16'h15a5] = 8'hca; ram[16'h15a6] = 8'hca; ram[16'h15a7] = 8'hca; 
ram[16'h15a8] = 8'hd0; ram[16'h15a9] = 8'hfe; ram[16'h15aa] = 8'ha9; ram[16'h15ab] = 8'h00; ram[16'h15ac] = 8'h48; ram[16'h15ad] = 8'ha9; ram[16'h15ae] = 8'h44; ram[16'h15af] = 8'h28; 
ram[16'h15b0] = 8'hbb; ram[16'h15b1] = 8'hea; ram[16'h15b2] = 8'hea; ram[16'h15b3] = 8'h08; ram[16'h15b4] = 8'hc9; ram[16'h15b5] = 8'h44; ram[16'h15b6] = 8'hd0; ram[16'h15b7] = 8'hfe; 
ram[16'h15b8] = 8'h68; ram[16'h15b9] = 8'h48; ram[16'h15ba] = 8'hc9; ram[16'h15bb] = 8'h30; ram[16'h15bc] = 8'hd0; ram[16'h15bd] = 8'hfe; ram[16'h15be] = 8'h28; ram[16'h15bf] = 8'ha9; 

ram[16'h15c0] = 8'hff; ram[16'h15c1] = 8'h48; ram[16'h15c2] = 8'ha9; ram[16'h15c3] = 8'hef; ram[16'h15c4] = 8'h28; ram[16'h15c5] = 8'hbb; ram[16'h15c6] = 8'hea; ram[16'h15c7] = 8'hea; 
ram[16'h15c8] = 8'h08; ram[16'h15c9] = 8'hc9; ram[16'h15ca] = 8'hef; ram[16'h15cb] = 8'hd0; ram[16'h15cc] = 8'hfe; ram[16'h15cd] = 8'h68; ram[16'h15ce] = 8'h48; ram[16'h15cf] = 8'hc9; 
ram[16'h15d0] = 8'hff; ram[16'h15d1] = 8'hd0; ram[16'h15d2] = 8'hfe; ram[16'h15d3] = 8'h28; ram[16'h15d4] = 8'hc0; ram[16'h15d5] = 8'h42; ram[16'h15d6] = 8'hd0; ram[16'h15d7] = 8'hfe; 
ram[16'h15d8] = 8'he0; ram[16'h15d9] = 8'h00; ram[16'h15da] = 8'hd0; ram[16'h15db] = 8'hfe; ram[16'h15dc] = 8'ha0; ram[16'h15dd] = 8'h42; ram[16'h15de] = 8'ha2; ram[16'h15df] = 8'h03; 

ram[16'h15e0] = 8'heb; ram[16'h15e1] = 8'hca; ram[16'h15e2] = 8'hca; ram[16'h15e3] = 8'hca; ram[16'h15e4] = 8'hd0; ram[16'h15e5] = 8'hfe; ram[16'h15e6] = 8'ha9; ram[16'h15e7] = 8'h00; 
ram[16'h15e8] = 8'h48; ram[16'h15e9] = 8'ha9; ram[16'h15ea] = 8'h14; ram[16'h15eb] = 8'h28; ram[16'h15ec] = 8'heb; ram[16'h15ed] = 8'hea; ram[16'h15ee] = 8'hea; ram[16'h15ef] = 8'h08; 
ram[16'h15f0] = 8'hc9; ram[16'h15f1] = 8'h14; ram[16'h15f2] = 8'hd0; ram[16'h15f3] = 8'hfe; ram[16'h15f4] = 8'h68; ram[16'h15f5] = 8'h48; ram[16'h15f6] = 8'hc9; ram[16'h15f7] = 8'h30; 
ram[16'h15f8] = 8'hd0; ram[16'h15f9] = 8'hfe; ram[16'h15fa] = 8'h28; ram[16'h15fb] = 8'ha9; ram[16'h15fc] = 8'hff; ram[16'h15fd] = 8'h48; ram[16'h15fe] = 8'ha9; ram[16'h15ff] = 8'hbf; 

ram[16'h1600] = 8'h28; ram[16'h1601] = 8'heb; ram[16'h1602] = 8'hea; ram[16'h1603] = 8'hea; ram[16'h1604] = 8'h08; ram[16'h1605] = 8'hc9; ram[16'h1606] = 8'hbf; ram[16'h1607] = 8'hd0; 
ram[16'h1608] = 8'hfe; ram[16'h1609] = 8'h68; ram[16'h160a] = 8'h48; ram[16'h160b] = 8'hc9; ram[16'h160c] = 8'hff; ram[16'h160d] = 8'hd0; ram[16'h160e] = 8'hfe; ram[16'h160f] = 8'h28; 
ram[16'h1610] = 8'hc0; ram[16'h1611] = 8'h42; ram[16'h1612] = 8'hd0; ram[16'h1613] = 8'hfe; ram[16'h1614] = 8'he0; ram[16'h1615] = 8'h00; ram[16'h1616] = 8'hd0; ram[16'h1617] = 8'hfe; 
ram[16'h1618] = 8'ha0; ram[16'h1619] = 8'h42; ram[16'h161a] = 8'ha2; ram[16'h161b] = 8'h03; ram[16'h161c] = 8'hfb; ram[16'h161d] = 8'hca; ram[16'h161e] = 8'hca; ram[16'h161f] = 8'hca; 

ram[16'h1620] = 8'hd0; ram[16'h1621] = 8'hfe; ram[16'h1622] = 8'ha9; ram[16'h1623] = 8'h00; ram[16'h1624] = 8'h48; ram[16'h1625] = 8'ha9; ram[16'h1626] = 8'h04; ram[16'h1627] = 8'h28; 
ram[16'h1628] = 8'hfb; ram[16'h1629] = 8'hea; ram[16'h162a] = 8'hea; ram[16'h162b] = 8'h08; ram[16'h162c] = 8'hc9; ram[16'h162d] = 8'h04; ram[16'h162e] = 8'hd0; ram[16'h162f] = 8'hfe; 
ram[16'h1630] = 8'h68; ram[16'h1631] = 8'h48; ram[16'h1632] = 8'hc9; ram[16'h1633] = 8'h30; ram[16'h1634] = 8'hd0; ram[16'h1635] = 8'hfe; ram[16'h1636] = 8'h28; ram[16'h1637] = 8'ha9; 
ram[16'h1638] = 8'hff; ram[16'h1639] = 8'h48; ram[16'h163a] = 8'ha9; ram[16'h163b] = 8'haf; ram[16'h163c] = 8'h28; ram[16'h163d] = 8'hfb; ram[16'h163e] = 8'hea; ram[16'h163f] = 8'hea; 

ram[16'h1640] = 8'h08; ram[16'h1641] = 8'hc9; ram[16'h1642] = 8'haf; ram[16'h1643] = 8'hd0; ram[16'h1644] = 8'hfe; ram[16'h1645] = 8'h68; ram[16'h1646] = 8'h48; ram[16'h1647] = 8'hc9; 
ram[16'h1648] = 8'hff; ram[16'h1649] = 8'hd0; ram[16'h164a] = 8'hfe; ram[16'h164b] = 8'h28; ram[16'h164c] = 8'hc0; ram[16'h164d] = 8'h42; ram[16'h164e] = 8'hd0; ram[16'h164f] = 8'hfe; 
ram[16'h1650] = 8'he0; ram[16'h1651] = 8'h00; ram[16'h1652] = 8'hd0; ram[16'h1653] = 8'hfe; ram[16'h1654] = 8'had; ram[16'h1655] = 8'h02; ram[16'h1656] = 8'h02; ram[16'h1657] = 8'hc9; 
ram[16'h1658] = 8'h08; ram[16'h1659] = 8'hd0; ram[16'h165a] = 8'hfe; ram[16'h165b] = 8'ha9; ram[16'h165c] = 8'h09; ram[16'h165d] = 8'h8d; ram[16'h165e] = 8'h02; ram[16'h165f] = 8'h02; 

ram[16'h1660] = 8'ha2; ram[16'h1661] = 8'h03; ram[16'h1662] = 8'hbd; ram[16'h1663] = 8'h8b; ram[16'h1664] = 8'h26; ram[16'h1665] = 8'h9d; ram[16'h1666] = 8'hfd; ram[16'h1667] = 8'h02; 
ram[16'h1668] = 8'hca; ram[16'h1669] = 8'h10; ram[16'h166a] = 8'hf7; ram[16'h166b] = 8'ha9; ram[16'h166c] = 8'h28; ram[16'h166d] = 8'h8d; ram[16'h166e] = 8'h00; ram[16'h166f] = 8'h02; 
ram[16'h1670] = 8'ha9; ram[16'h1671] = 8'h00; ram[16'h1672] = 8'h48; ram[16'h1673] = 8'h28; ram[16'h1674] = 8'ha9; ram[16'h1675] = 8'h49; ram[16'h1676] = 8'ha2; ram[16'h1677] = 8'h4e; 
ram[16'h1678] = 8'ha0; ram[16'h1679] = 8'h44; ram[16'h167a] = 8'h6c; ram[16'h167b] = 8'hfd; ram[16'h167c] = 8'h02; ram[16'h167d] = 8'hea; ram[16'h167e] = 8'hd0; ram[16'h167f] = 8'hfe; 

ram[16'h1680] = 8'h88; ram[16'h1681] = 8'h88; ram[16'h1682] = 8'h08; ram[16'h1683] = 8'h88; ram[16'h1684] = 8'h88; ram[16'h1685] = 8'h88; ram[16'h1686] = 8'h28; ram[16'h1687] = 8'hf0; 
ram[16'h1688] = 8'hfe; ram[16'h1689] = 8'h10; ram[16'h168a] = 8'hfe; ram[16'h168b] = 8'h90; ram[16'h168c] = 8'hfe; ram[16'h168d] = 8'h50; ram[16'h168e] = 8'hfe; ram[16'h168f] = 8'hc9; 
ram[16'h1690] = 8'he3; ram[16'h1691] = 8'hd0; ram[16'h1692] = 8'hfe; ram[16'h1693] = 8'he0; ram[16'h1694] = 8'h4f; ram[16'h1695] = 8'hd0; ram[16'h1696] = 8'hfe; ram[16'h1697] = 8'hc0; 
ram[16'h1698] = 8'h3e; ram[16'h1699] = 8'hd0; ram[16'h169a] = 8'hfe; ram[16'h169b] = 8'hba; ram[16'h169c] = 8'he0; ram[16'h169d] = 8'hff; ram[16'h169e] = 8'hd0; ram[16'h169f] = 8'hfe; 

ram[16'h16a0] = 8'had; ram[16'h16a1] = 8'h02; ram[16'h16a2] = 8'h02; ram[16'h16a3] = 8'hc9; ram[16'h16a4] = 8'h09; ram[16'h16a5] = 8'hd0; ram[16'h16a6] = 8'hfe; ram[16'h16a7] = 8'ha9; 
ram[16'h16a8] = 8'h0a; ram[16'h16a9] = 8'h8d; ram[16'h16aa] = 8'h02; ram[16'h16ab] = 8'h02; ram[16'h16ac] = 8'ha2; ram[16'h16ad] = 8'h0b; ram[16'h16ae] = 8'hbd; ram[16'h16af] = 8'hc7; 
ram[16'h16b0] = 8'h26; ram[16'h16b1] = 8'h9d; ram[16'h16b2] = 8'hf9; ram[16'h16b3] = 8'h02; ram[16'h16b4] = 8'hca; ram[16'h16b5] = 8'h10; ram[16'h16b6] = 8'hf7; ram[16'h16b7] = 8'ha9; 
ram[16'h16b8] = 8'h27; ram[16'h16b9] = 8'h8d; ram[16'h16ba] = 8'h00; ram[16'h16bb] = 8'h02; ram[16'h16bc] = 8'ha9; ram[16'h16bd] = 8'h00; ram[16'h16be] = 8'h48; ram[16'h16bf] = 8'h28; 

ram[16'h16c0] = 8'ha9; ram[16'h16c1] = 8'h58; ram[16'h16c2] = 8'ha2; ram[16'h16c3] = 8'h04; ram[16'h16c4] = 8'ha0; ram[16'h16c5] = 8'h49; ram[16'h16c6] = 8'h7c; ram[16'h16c7] = 8'hf9; 
ram[16'h16c8] = 8'h02; ram[16'h16c9] = 8'hea; ram[16'h16ca] = 8'hd0; ram[16'h16cb] = 8'hfe; ram[16'h16cc] = 8'h88; ram[16'h16cd] = 8'h88; ram[16'h16ce] = 8'h08; ram[16'h16cf] = 8'h88; 
ram[16'h16d0] = 8'h88; ram[16'h16d1] = 8'h88; ram[16'h16d2] = 8'h28; ram[16'h16d3] = 8'hf0; ram[16'h16d4] = 8'hfe; ram[16'h16d5] = 8'h10; ram[16'h16d6] = 8'hfe; ram[16'h16d7] = 8'h90; 
ram[16'h16d8] = 8'hfe; ram[16'h16d9] = 8'h50; ram[16'h16da] = 8'hfe; ram[16'h16db] = 8'hc9; ram[16'h16dc] = 8'hf2; ram[16'h16dd] = 8'hd0; ram[16'h16de] = 8'hfe; ram[16'h16df] = 8'he0; 

ram[16'h16e0] = 8'h06; ram[16'h16e1] = 8'hd0; ram[16'h16e2] = 8'hfe; ram[16'h16e3] = 8'hc0; ram[16'h16e4] = 8'h43; ram[16'h16e5] = 8'hd0; ram[16'h16e6] = 8'hfe; ram[16'h16e7] = 8'hba; 
ram[16'h16e8] = 8'he0; ram[16'h16e9] = 8'hff; ram[16'h16ea] = 8'hd0; ram[16'h16eb] = 8'hfe; ram[16'h16ec] = 8'ha9; ram[16'h16ed] = 8'h08; ram[16'h16ee] = 8'h8d; ram[16'h16ef] = 8'h00; 
ram[16'h16f0] = 8'h03; ram[16'h16f1] = 8'ha9; ram[16'h16f2] = 8'h17; ram[16'h16f3] = 8'h8d; ram[16'h16f4] = 8'h01; ram[16'h16f5] = 8'h03; ram[16'h16f6] = 8'ha9; ram[16'h16f7] = 8'h05; 
ram[16'h16f8] = 8'h8d; ram[16'h16f9] = 8'h00; ram[16'h16fa] = 8'h02; ram[16'h16fb] = 8'ha9; ram[16'h16fc] = 8'h17; ram[16'h16fd] = 8'h8d; ram[16'h16fe] = 8'h01; ram[16'h16ff] = 8'h02; 

ram[16'h1700] = 8'ha2; ram[16'h1701] = 8'hff; ram[16'h1702] = 8'h7c; ram[16'h1703] = 8'h01; ram[16'h1704] = 8'h02; ram[16'h1705] = 8'h4c; ram[16'h1706] = 8'h05; ram[16'h1707] = 8'h17; 
ram[16'h1708] = 8'had; ram[16'h1709] = 8'h02; ram[16'h170a] = 8'h02; ram[16'h170b] = 8'hc9; ram[16'h170c] = 8'h0a; ram[16'h170d] = 8'hd0; ram[16'h170e] = 8'hfe; ram[16'h170f] = 8'ha9; 
ram[16'h1710] = 8'h0b; ram[16'h1711] = 8'h8d; ram[16'h1712] = 8'h02; ram[16'h1713] = 8'h02; ram[16'h1714] = 8'ha9; ram[16'h1715] = 8'h00; ram[16'h1716] = 8'h48; ram[16'h1717] = 8'ha9; 
ram[16'h1718] = 8'h42; ram[16'h1719] = 8'ha2; ram[16'h171a] = 8'h52; ram[16'h171b] = 8'ha0; ram[16'h171c] = 8'h4b; ram[16'h171d] = 8'h28; ram[16'h171e] = 8'h00; ram[16'h171f] = 8'h88; 

ram[16'h1720] = 8'h08; ram[16'h1721] = 8'h88; ram[16'h1722] = 8'h88; ram[16'h1723] = 8'h88; ram[16'h1724] = 8'hc9; ram[16'h1725] = 8'he8; ram[16'h1726] = 8'hd0; ram[16'h1727] = 8'hfe; 
ram[16'h1728] = 8'he0; ram[16'h1729] = 8'h53; ram[16'h172a] = 8'hd0; ram[16'h172b] = 8'hfe; ram[16'h172c] = 8'hc0; ram[16'h172d] = 8'h45; ram[16'h172e] = 8'hd0; ram[16'h172f] = 8'hfe; 
ram[16'h1730] = 8'h68; ram[16'h1731] = 8'hc9; ram[16'h1732] = 8'h30; ram[16'h1733] = 8'hd0; ram[16'h1734] = 8'hfe; ram[16'h1735] = 8'hba; ram[16'h1736] = 8'he0; ram[16'h1737] = 8'hff; 
ram[16'h1738] = 8'hd0; ram[16'h1739] = 8'hfe; ram[16'h173a] = 8'ha9; ram[16'h173b] = 8'hff; ram[16'h173c] = 8'h48; ram[16'h173d] = 8'ha9; ram[16'h173e] = 8'hbd; ram[16'h173f] = 8'ha2; 

ram[16'h1740] = 8'had; ram[16'h1741] = 8'ha0; ram[16'h1742] = 8'hb4; ram[16'h1743] = 8'h28; ram[16'h1744] = 8'h00; ram[16'h1745] = 8'h88; ram[16'h1746] = 8'h08; ram[16'h1747] = 8'h88; 
ram[16'h1748] = 8'h88; ram[16'h1749] = 8'h88; ram[16'h174a] = 8'hc9; ram[16'h174b] = 8'h17; ram[16'h174c] = 8'hd0; ram[16'h174d] = 8'hfe; ram[16'h174e] = 8'he0; ram[16'h174f] = 8'hae; 
ram[16'h1750] = 8'hd0; ram[16'h1751] = 8'hfe; ram[16'h1752] = 8'hc0; ram[16'h1753] = 8'hae; ram[16'h1754] = 8'hd0; ram[16'h1755] = 8'hfe; ram[16'h1756] = 8'h68; ram[16'h1757] = 8'hc9; 
ram[16'h1758] = 8'hff; ram[16'h1759] = 8'hd0; ram[16'h175a] = 8'hfe; ram[16'h175b] = 8'hba; ram[16'h175c] = 8'he0; ram[16'h175d] = 8'hff; ram[16'h175e] = 8'hd0; ram[16'h175f] = 8'hfe; 

ram[16'h1760] = 8'had; ram[16'h1761] = 8'h02; ram[16'h1762] = 8'h02; ram[16'h1763] = 8'hc9; ram[16'h1764] = 8'h0b; ram[16'h1765] = 8'hd0; ram[16'h1766] = 8'hfe; ram[16'h1767] = 8'ha9; 
ram[16'h1768] = 8'h0c; ram[16'h1769] = 8'h8d; ram[16'h176a] = 8'h02; ram[16'h176b] = 8'h02; ram[16'h176c] = 8'ha2; ram[16'h176d] = 8'hac; ram[16'h176e] = 8'ha0; ram[16'h176f] = 8'hdc; 
ram[16'h1770] = 8'ha9; ram[16'h1771] = 8'hff; ram[16'h1772] = 8'h48; ram[16'h1773] = 8'ha9; ram[16'h1774] = 8'hfe; ram[16'h1775] = 8'h28; ram[16'h1776] = 8'h1a; ram[16'h1777] = 8'h48; 
ram[16'h1778] = 8'h08; ram[16'h1779] = 8'hc9; ram[16'h177a] = 8'hff; ram[16'h177b] = 8'hd0; ram[16'h177c] = 8'hfe; ram[16'h177d] = 8'h68; ram[16'h177e] = 8'h48; ram[16'h177f] = 8'hc9; 

ram[16'h1780] = 8'hfd; ram[16'h1781] = 8'hd0; ram[16'h1782] = 8'hfe; ram[16'h1783] = 8'h28; ram[16'h1784] = 8'h68; ram[16'h1785] = 8'h1a; ram[16'h1786] = 8'h48; ram[16'h1787] = 8'h08; 
ram[16'h1788] = 8'hc9; ram[16'h1789] = 8'h00; ram[16'h178a] = 8'hd0; ram[16'h178b] = 8'hfe; ram[16'h178c] = 8'h68; ram[16'h178d] = 8'h48; ram[16'h178e] = 8'hc9; ram[16'h178f] = 8'h7f; 
ram[16'h1790] = 8'hd0; ram[16'h1791] = 8'hfe; ram[16'h1792] = 8'h28; ram[16'h1793] = 8'h68; ram[16'h1794] = 8'h1a; ram[16'h1795] = 8'h48; ram[16'h1796] = 8'h08; ram[16'h1797] = 8'hc9; 
ram[16'h1798] = 8'h01; ram[16'h1799] = 8'hd0; ram[16'h179a] = 8'hfe; ram[16'h179b] = 8'h68; ram[16'h179c] = 8'h48; ram[16'h179d] = 8'hc9; ram[16'h179e] = 8'h7d; ram[16'h179f] = 8'hd0; 

ram[16'h17a0] = 8'hfe; ram[16'h17a1] = 8'h28; ram[16'h17a2] = 8'h68; ram[16'h17a3] = 8'h3a; ram[16'h17a4] = 8'h48; ram[16'h17a5] = 8'h08; ram[16'h17a6] = 8'hc9; ram[16'h17a7] = 8'h00; 
ram[16'h17a8] = 8'hd0; ram[16'h17a9] = 8'hfe; ram[16'h17aa] = 8'h68; ram[16'h17ab] = 8'h48; ram[16'h17ac] = 8'hc9; ram[16'h17ad] = 8'h7f; ram[16'h17ae] = 8'hd0; ram[16'h17af] = 8'hfe; 
ram[16'h17b0] = 8'h28; ram[16'h17b1] = 8'h68; ram[16'h17b2] = 8'h3a; ram[16'h17b3] = 8'h48; ram[16'h17b4] = 8'h08; ram[16'h17b5] = 8'hc9; ram[16'h17b6] = 8'hff; ram[16'h17b7] = 8'hd0; 
ram[16'h17b8] = 8'hfe; ram[16'h17b9] = 8'h68; ram[16'h17ba] = 8'h48; ram[16'h17bb] = 8'hc9; ram[16'h17bc] = 8'hfd; ram[16'h17bd] = 8'hd0; ram[16'h17be] = 8'hfe; ram[16'h17bf] = 8'h28; 

ram[16'h17c0] = 8'h68; ram[16'h17c1] = 8'h3a; ram[16'h17c2] = 8'ha9; ram[16'h17c3] = 8'h00; ram[16'h17c4] = 8'h48; ram[16'h17c5] = 8'ha9; ram[16'h17c6] = 8'hfe; ram[16'h17c7] = 8'h28; 
ram[16'h17c8] = 8'h1a; ram[16'h17c9] = 8'h48; ram[16'h17ca] = 8'h08; ram[16'h17cb] = 8'hc9; ram[16'h17cc] = 8'hff; ram[16'h17cd] = 8'hd0; ram[16'h17ce] = 8'hfe; ram[16'h17cf] = 8'h68; 
ram[16'h17d0] = 8'h48; ram[16'h17d1] = 8'hc9; ram[16'h17d2] = 8'hb0; ram[16'h17d3] = 8'hd0; ram[16'h17d4] = 8'hfe; ram[16'h17d5] = 8'h28; ram[16'h17d6] = 8'h68; ram[16'h17d7] = 8'h1a; 
ram[16'h17d8] = 8'h48; ram[16'h17d9] = 8'h08; ram[16'h17da] = 8'hc9; ram[16'h17db] = 8'h00; ram[16'h17dc] = 8'hd0; ram[16'h17dd] = 8'hfe; ram[16'h17de] = 8'h68; ram[16'h17df] = 8'h48; 

ram[16'h17e0] = 8'hc9; ram[16'h17e1] = 8'h32; ram[16'h17e2] = 8'hd0; ram[16'h17e3] = 8'hfe; ram[16'h17e4] = 8'h28; ram[16'h17e5] = 8'h68; ram[16'h17e6] = 8'h1a; ram[16'h17e7] = 8'h48; 
ram[16'h17e8] = 8'h08; ram[16'h17e9] = 8'hc9; ram[16'h17ea] = 8'h01; ram[16'h17eb] = 8'hd0; ram[16'h17ec] = 8'hfe; ram[16'h17ed] = 8'h68; ram[16'h17ee] = 8'h48; ram[16'h17ef] = 8'hc9; 
ram[16'h17f0] = 8'h30; ram[16'h17f1] = 8'hd0; ram[16'h17f2] = 8'hfe; ram[16'h17f3] = 8'h28; ram[16'h17f4] = 8'h68; ram[16'h17f5] = 8'h3a; ram[16'h17f6] = 8'h48; ram[16'h17f7] = 8'h08; 
ram[16'h17f8] = 8'hc9; ram[16'h17f9] = 8'h00; ram[16'h17fa] = 8'hd0; ram[16'h17fb] = 8'hfe; ram[16'h17fc] = 8'h68; ram[16'h17fd] = 8'h48; ram[16'h17fe] = 8'hc9; ram[16'h17ff] = 8'h32; 

ram[16'h1800] = 8'hd0; ram[16'h1801] = 8'hfe; ram[16'h1802] = 8'h28; ram[16'h1803] = 8'h68; ram[16'h1804] = 8'h3a; ram[16'h1805] = 8'h48; ram[16'h1806] = 8'h08; ram[16'h1807] = 8'hc9; 
ram[16'h1808] = 8'hff; ram[16'h1809] = 8'hd0; ram[16'h180a] = 8'hfe; ram[16'h180b] = 8'h68; ram[16'h180c] = 8'h48; ram[16'h180d] = 8'hc9; ram[16'h180e] = 8'hb0; ram[16'h180f] = 8'hd0; 
ram[16'h1810] = 8'hfe; ram[16'h1811] = 8'h28; ram[16'h1812] = 8'h68; ram[16'h1813] = 8'he0; ram[16'h1814] = 8'hac; ram[16'h1815] = 8'hd0; ram[16'h1816] = 8'hfe; ram[16'h1817] = 8'hc0; 
ram[16'h1818] = 8'hdc; ram[16'h1819] = 8'hd0; ram[16'h181a] = 8'hfe; ram[16'h181b] = 8'hba; ram[16'h181c] = 8'he0; ram[16'h181d] = 8'hff; ram[16'h181e] = 8'hd0; ram[16'h181f] = 8'hfe; 

ram[16'h1820] = 8'had; ram[16'h1821] = 8'h02; ram[16'h1822] = 8'h02; ram[16'h1823] = 8'hc9; ram[16'h1824] = 8'h0c; ram[16'h1825] = 8'hd0; ram[16'h1826] = 8'hfe; ram[16'h1827] = 8'ha9; 
ram[16'h1828] = 8'h0d; ram[16'h1829] = 8'h8d; ram[16'h182a] = 8'h02; ram[16'h182b] = 8'h02; ram[16'h182c] = 8'ha2; ram[16'h182d] = 8'h99; ram[16'h182e] = 8'ha0; ram[16'h182f] = 8'h66; 
ram[16'h1830] = 8'ha9; ram[16'h1831] = 8'h00; ram[16'h1832] = 8'h48; ram[16'h1833] = 8'h28; ram[16'h1834] = 8'hb2; ram[16'h1835] = 8'h24; ram[16'h1836] = 8'h08; ram[16'h1837] = 8'h49; 
ram[16'h1838] = 8'hc3; ram[16'h1839] = 8'h28; ram[16'h183a] = 8'h92; ram[16'h183b] = 8'h30; ram[16'h183c] = 8'h08; ram[16'h183d] = 8'h49; ram[16'h183e] = 8'hc3; ram[16'h183f] = 8'hc9; 

ram[16'h1840] = 8'hc3; ram[16'h1841] = 8'hd0; ram[16'h1842] = 8'hfe; ram[16'h1843] = 8'h68; ram[16'h1844] = 8'h49; ram[16'h1845] = 8'h30; ram[16'h1846] = 8'hcd; ram[16'h1847] = 8'h15; 
ram[16'h1848] = 8'h02; ram[16'h1849] = 8'hd0; ram[16'h184a] = 8'hfe; ram[16'h184b] = 8'ha9; ram[16'h184c] = 8'h00; ram[16'h184d] = 8'h48; ram[16'h184e] = 8'h28; ram[16'h184f] = 8'hb2; 
ram[16'h1850] = 8'h26; ram[16'h1851] = 8'h08; ram[16'h1852] = 8'h49; ram[16'h1853] = 8'hc3; ram[16'h1854] = 8'h28; ram[16'h1855] = 8'h92; ram[16'h1856] = 8'h32; ram[16'h1857] = 8'h08; 
ram[16'h1858] = 8'h49; ram[16'h1859] = 8'hc3; ram[16'h185a] = 8'hc9; ram[16'h185b] = 8'h82; ram[16'h185c] = 8'hd0; ram[16'h185d] = 8'hfe; ram[16'h185e] = 8'h68; ram[16'h185f] = 8'h49; 

ram[16'h1860] = 8'h30; ram[16'h1861] = 8'hcd; ram[16'h1862] = 8'h16; ram[16'h1863] = 8'h02; ram[16'h1864] = 8'hd0; ram[16'h1865] = 8'hfe; ram[16'h1866] = 8'ha9; ram[16'h1867] = 8'h00; 
ram[16'h1868] = 8'h48; ram[16'h1869] = 8'h28; ram[16'h186a] = 8'hb2; ram[16'h186b] = 8'h28; ram[16'h186c] = 8'h08; ram[16'h186d] = 8'h49; ram[16'h186e] = 8'hc3; ram[16'h186f] = 8'h28; 
ram[16'h1870] = 8'h92; ram[16'h1871] = 8'h34; ram[16'h1872] = 8'h08; ram[16'h1873] = 8'h49; ram[16'h1874] = 8'hc3; ram[16'h1875] = 8'hc9; ram[16'h1876] = 8'h41; ram[16'h1877] = 8'hd0; 
ram[16'h1878] = 8'hfe; ram[16'h1879] = 8'h68; ram[16'h187a] = 8'h49; ram[16'h187b] = 8'h30; ram[16'h187c] = 8'hcd; ram[16'h187d] = 8'h17; ram[16'h187e] = 8'h02; ram[16'h187f] = 8'hd0; 

ram[16'h1880] = 8'hfe; ram[16'h1881] = 8'ha9; ram[16'h1882] = 8'h00; ram[16'h1883] = 8'h48; ram[16'h1884] = 8'h28; ram[16'h1885] = 8'hb2; ram[16'h1886] = 8'h2a; ram[16'h1887] = 8'h08; 
ram[16'h1888] = 8'h49; ram[16'h1889] = 8'hc3; ram[16'h188a] = 8'h28; ram[16'h188b] = 8'h92; ram[16'h188c] = 8'h36; ram[16'h188d] = 8'h08; ram[16'h188e] = 8'h49; ram[16'h188f] = 8'hc3; 
ram[16'h1890] = 8'hc9; ram[16'h1891] = 8'h00; ram[16'h1892] = 8'hd0; ram[16'h1893] = 8'hfe; ram[16'h1894] = 8'h68; ram[16'h1895] = 8'h49; ram[16'h1896] = 8'h30; ram[16'h1897] = 8'hcd; 
ram[16'h1898] = 8'h18; ram[16'h1899] = 8'h02; ram[16'h189a] = 8'hd0; ram[16'h189b] = 8'hfe; ram[16'h189c] = 8'he0; ram[16'h189d] = 8'h99; ram[16'h189e] = 8'hd0; ram[16'h189f] = 8'hfe; 

ram[16'h18a0] = 8'hc0; ram[16'h18a1] = 8'h66; ram[16'h18a2] = 8'hd0; ram[16'h18a3] = 8'hfe; ram[16'h18a4] = 8'ha0; ram[16'h18a5] = 8'h03; ram[16'h18a6] = 8'ha2; ram[16'h18a7] = 8'h00; 
ram[16'h18a8] = 8'hb9; ram[16'h18a9] = 8'h05; ram[16'h18aa] = 8'h02; ram[16'h18ab] = 8'h49; ram[16'h18ac] = 8'hc3; ram[16'h18ad] = 8'hd9; ram[16'h18ae] = 8'h10; ram[16'h18af] = 8'h02; 
ram[16'h18b0] = 8'hd0; ram[16'h18b1] = 8'hfe; ram[16'h18b2] = 8'h8a; ram[16'h18b3] = 8'h99; ram[16'h18b4] = 8'h05; ram[16'h18b5] = 8'h02; ram[16'h18b6] = 8'h88; ram[16'h18b7] = 8'h10; 
ram[16'h18b8] = 8'hef; ram[16'h18b9] = 8'ha2; ram[16'h18ba] = 8'h99; ram[16'h18bb] = 8'ha0; ram[16'h18bc] = 8'h66; ram[16'h18bd] = 8'ha9; ram[16'h18be] = 8'hff; ram[16'h18bf] = 8'h48; 

ram[16'h18c0] = 8'h28; ram[16'h18c1] = 8'hb2; ram[16'h18c2] = 8'h24; ram[16'h18c3] = 8'h08; ram[16'h18c4] = 8'h49; ram[16'h18c5] = 8'hc3; ram[16'h18c6] = 8'h28; ram[16'h18c7] = 8'h92; 
ram[16'h18c8] = 8'h30; ram[16'h18c9] = 8'h08; ram[16'h18ca] = 8'h49; ram[16'h18cb] = 8'hc3; ram[16'h18cc] = 8'hc9; ram[16'h18cd] = 8'hc3; ram[16'h18ce] = 8'hd0; ram[16'h18cf] = 8'hfe; 
ram[16'h18d0] = 8'h68; ram[16'h18d1] = 8'h49; ram[16'h18d2] = 8'h7d; ram[16'h18d3] = 8'hcd; ram[16'h18d4] = 8'h15; ram[16'h18d5] = 8'h02; ram[16'h18d6] = 8'hd0; ram[16'h18d7] = 8'hfe; 
ram[16'h18d8] = 8'ha9; ram[16'h18d9] = 8'hff; ram[16'h18da] = 8'h48; ram[16'h18db] = 8'h28; ram[16'h18dc] = 8'hb2; ram[16'h18dd] = 8'h26; ram[16'h18de] = 8'h08; ram[16'h18df] = 8'h49; 

ram[16'h18e0] = 8'hc3; ram[16'h18e1] = 8'h28; ram[16'h18e2] = 8'h92; ram[16'h18e3] = 8'h32; ram[16'h18e4] = 8'h08; ram[16'h18e5] = 8'h49; ram[16'h18e6] = 8'hc3; ram[16'h18e7] = 8'hc9; 
ram[16'h18e8] = 8'h82; ram[16'h18e9] = 8'hd0; ram[16'h18ea] = 8'hfe; ram[16'h18eb] = 8'h68; ram[16'h18ec] = 8'h49; ram[16'h18ed] = 8'h7d; ram[16'h18ee] = 8'hcd; ram[16'h18ef] = 8'h16; 
ram[16'h18f0] = 8'h02; ram[16'h18f1] = 8'hd0; ram[16'h18f2] = 8'hfe; ram[16'h18f3] = 8'ha9; ram[16'h18f4] = 8'hff; ram[16'h18f5] = 8'h48; ram[16'h18f6] = 8'h28; ram[16'h18f7] = 8'hb2; 
ram[16'h18f8] = 8'h28; ram[16'h18f9] = 8'h08; ram[16'h18fa] = 8'h49; ram[16'h18fb] = 8'hc3; ram[16'h18fc] = 8'h28; ram[16'h18fd] = 8'h92; ram[16'h18fe] = 8'h34; ram[16'h18ff] = 8'h08; 

ram[16'h1900] = 8'h49; ram[16'h1901] = 8'hc3; ram[16'h1902] = 8'hc9; ram[16'h1903] = 8'h41; ram[16'h1904] = 8'hd0; ram[16'h1905] = 8'hfe; ram[16'h1906] = 8'h68; ram[16'h1907] = 8'h49; 
ram[16'h1908] = 8'h7d; ram[16'h1909] = 8'hcd; ram[16'h190a] = 8'h17; ram[16'h190b] = 8'h02; ram[16'h190c] = 8'hd0; ram[16'h190d] = 8'hfe; ram[16'h190e] = 8'ha9; ram[16'h190f] = 8'hff; 
ram[16'h1910] = 8'h48; ram[16'h1911] = 8'h28; ram[16'h1912] = 8'hb2; ram[16'h1913] = 8'h2a; ram[16'h1914] = 8'h08; ram[16'h1915] = 8'h49; ram[16'h1916] = 8'hc3; ram[16'h1917] = 8'h28; 
ram[16'h1918] = 8'h92; ram[16'h1919] = 8'h36; ram[16'h191a] = 8'h08; ram[16'h191b] = 8'h49; ram[16'h191c] = 8'hc3; ram[16'h191d] = 8'hc9; ram[16'h191e] = 8'h00; ram[16'h191f] = 8'hd0; 

ram[16'h1920] = 8'hfe; ram[16'h1921] = 8'h68; ram[16'h1922] = 8'h49; ram[16'h1923] = 8'h7d; ram[16'h1924] = 8'hcd; ram[16'h1925] = 8'h18; ram[16'h1926] = 8'h02; ram[16'h1927] = 8'hd0; 
ram[16'h1928] = 8'hfe; ram[16'h1929] = 8'he0; ram[16'h192a] = 8'h99; ram[16'h192b] = 8'hd0; ram[16'h192c] = 8'hfe; ram[16'h192d] = 8'hc0; ram[16'h192e] = 8'h66; ram[16'h192f] = 8'hd0; 
ram[16'h1930] = 8'hfe; ram[16'h1931] = 8'ha0; ram[16'h1932] = 8'h03; ram[16'h1933] = 8'ha2; ram[16'h1934] = 8'h00; ram[16'h1935] = 8'hb9; ram[16'h1936] = 8'h05; ram[16'h1937] = 8'h02; 
ram[16'h1938] = 8'h49; ram[16'h1939] = 8'hc3; ram[16'h193a] = 8'hd9; ram[16'h193b] = 8'h10; ram[16'h193c] = 8'h02; ram[16'h193d] = 8'hd0; ram[16'h193e] = 8'hfe; ram[16'h193f] = 8'h8a; 

ram[16'h1940] = 8'h99; ram[16'h1941] = 8'h05; ram[16'h1942] = 8'h02; ram[16'h1943] = 8'h88; ram[16'h1944] = 8'h10; ram[16'h1945] = 8'hef; ram[16'h1946] = 8'hba; ram[16'h1947] = 8'he0; 
ram[16'h1948] = 8'hff; ram[16'h1949] = 8'hd0; ram[16'h194a] = 8'hfe; ram[16'h194b] = 8'had; ram[16'h194c] = 8'h02; ram[16'h194d] = 8'h02; ram[16'h194e] = 8'hc9; ram[16'h194f] = 8'h0d; 
ram[16'h1950] = 8'hd0; ram[16'h1951] = 8'hfe; ram[16'h1952] = 8'ha9; ram[16'h1953] = 8'h0e; ram[16'h1954] = 8'h8d; ram[16'h1955] = 8'h02; ram[16'h1956] = 8'h02; ram[16'h1957] = 8'ha0; 
ram[16'h1958] = 8'h7b; ram[16'h1959] = 8'ha2; ram[16'h195a] = 8'h04; ram[16'h195b] = 8'ha9; ram[16'h195c] = 8'h07; ram[16'h195d] = 8'h95; ram[16'h195e] = 8'h0c; ram[16'h195f] = 8'h0a; 

ram[16'h1960] = 8'hca; ram[16'h1961] = 8'h10; ram[16'h1962] = 8'hfa; ram[16'h1963] = 8'ha2; ram[16'h1964] = 8'h04; ram[16'h1965] = 8'ha9; ram[16'h1966] = 8'hff; ram[16'h1967] = 8'h48; 
ram[16'h1968] = 8'ha9; ram[16'h1969] = 8'h55; ram[16'h196a] = 8'h28; ram[16'h196b] = 8'h64; ram[16'h196c] = 8'h0c; ram[16'h196d] = 8'h64; ram[16'h196e] = 8'h0d; ram[16'h196f] = 8'h64; 
ram[16'h1970] = 8'h0e; ram[16'h1971] = 8'h64; ram[16'h1972] = 8'h0f; ram[16'h1973] = 8'h64; ram[16'h1974] = 8'h10; ram[16'h1975] = 8'h08; ram[16'h1976] = 8'hc9; ram[16'h1977] = 8'h55; 
ram[16'h1978] = 8'hd0; ram[16'h1979] = 8'hfe; ram[16'h197a] = 8'h68; ram[16'h197b] = 8'h48; ram[16'h197c] = 8'hc9; ram[16'h197d] = 8'hff; ram[16'h197e] = 8'hd0; ram[16'h197f] = 8'hfe; 

ram[16'h1980] = 8'h28; ram[16'h1981] = 8'hb5; ram[16'h1982] = 8'h0c; ram[16'h1983] = 8'hd0; ram[16'h1984] = 8'hfe; ram[16'h1985] = 8'hca; ram[16'h1986] = 8'h10; ram[16'h1987] = 8'hf9; 
ram[16'h1988] = 8'ha2; ram[16'h1989] = 8'h04; ram[16'h198a] = 8'ha9; ram[16'h198b] = 8'h07; ram[16'h198c] = 8'h95; ram[16'h198d] = 8'h0c; ram[16'h198e] = 8'h0a; ram[16'h198f] = 8'hca; 
ram[16'h1990] = 8'h10; ram[16'h1991] = 8'hfa; ram[16'h1992] = 8'ha2; ram[16'h1993] = 8'h04; ram[16'h1994] = 8'ha9; ram[16'h1995] = 8'h00; ram[16'h1996] = 8'h48; ram[16'h1997] = 8'ha9; 
ram[16'h1998] = 8'haa; ram[16'h1999] = 8'h28; ram[16'h199a] = 8'h64; ram[16'h199b] = 8'h0c; ram[16'h199c] = 8'h64; ram[16'h199d] = 8'h0d; ram[16'h199e] = 8'h64; ram[16'h199f] = 8'h0e; 

ram[16'h19a0] = 8'h64; ram[16'h19a1] = 8'h0f; ram[16'h19a2] = 8'h64; ram[16'h19a3] = 8'h10; ram[16'h19a4] = 8'h08; ram[16'h19a5] = 8'hc9; ram[16'h19a6] = 8'haa; ram[16'h19a7] = 8'hd0; 
ram[16'h19a8] = 8'hfe; ram[16'h19a9] = 8'h68; ram[16'h19aa] = 8'h48; ram[16'h19ab] = 8'hc9; ram[16'h19ac] = 8'h30; ram[16'h19ad] = 8'hd0; ram[16'h19ae] = 8'hfe; ram[16'h19af] = 8'h28; 
ram[16'h19b0] = 8'hb5; ram[16'h19b1] = 8'h0c; ram[16'h19b2] = 8'hd0; ram[16'h19b3] = 8'hfe; ram[16'h19b4] = 8'hca; ram[16'h19b5] = 8'h10; ram[16'h19b6] = 8'hf9; ram[16'h19b7] = 8'ha2; 
ram[16'h19b8] = 8'h04; ram[16'h19b9] = 8'ha9; ram[16'h19ba] = 8'h07; ram[16'h19bb] = 8'h9d; ram[16'h19bc] = 8'h05; ram[16'h19bd] = 8'h02; ram[16'h19be] = 8'h0a; ram[16'h19bf] = 8'hca; 

ram[16'h19c0] = 8'h10; ram[16'h19c1] = 8'hf9; ram[16'h19c2] = 8'ha2; ram[16'h19c3] = 8'h04; ram[16'h19c4] = 8'ha9; ram[16'h19c5] = 8'hff; ram[16'h19c6] = 8'h48; ram[16'h19c7] = 8'ha9; 
ram[16'h19c8] = 8'h55; ram[16'h19c9] = 8'h28; ram[16'h19ca] = 8'h9c; ram[16'h19cb] = 8'h05; ram[16'h19cc] = 8'h02; ram[16'h19cd] = 8'h9c; ram[16'h19ce] = 8'h06; ram[16'h19cf] = 8'h02; 
ram[16'h19d0] = 8'h9c; ram[16'h19d1] = 8'h07; ram[16'h19d2] = 8'h02; ram[16'h19d3] = 8'h9c; ram[16'h19d4] = 8'h08; ram[16'h19d5] = 8'h02; ram[16'h19d6] = 8'h9c; ram[16'h19d7] = 8'h09; 
ram[16'h19d8] = 8'h02; ram[16'h19d9] = 8'h08; ram[16'h19da] = 8'hc9; ram[16'h19db] = 8'h55; ram[16'h19dc] = 8'hd0; ram[16'h19dd] = 8'hfe; ram[16'h19de] = 8'h68; ram[16'h19df] = 8'h48; 

ram[16'h19e0] = 8'hc9; ram[16'h19e1] = 8'hff; ram[16'h19e2] = 8'hd0; ram[16'h19e3] = 8'hfe; ram[16'h19e4] = 8'h28; ram[16'h19e5] = 8'hbd; ram[16'h19e6] = 8'h05; ram[16'h19e7] = 8'h02; 
ram[16'h19e8] = 8'hd0; ram[16'h19e9] = 8'hfe; ram[16'h19ea] = 8'hca; ram[16'h19eb] = 8'h10; ram[16'h19ec] = 8'hf8; ram[16'h19ed] = 8'ha2; ram[16'h19ee] = 8'h04; ram[16'h19ef] = 8'ha9; 
ram[16'h19f0] = 8'h07; ram[16'h19f1] = 8'h9d; ram[16'h19f2] = 8'h05; ram[16'h19f3] = 8'h02; ram[16'h19f4] = 8'h0a; ram[16'h19f5] = 8'hca; ram[16'h19f6] = 8'h10; ram[16'h19f7] = 8'hf9; 
ram[16'h19f8] = 8'ha2; ram[16'h19f9] = 8'h04; ram[16'h19fa] = 8'ha9; ram[16'h19fb] = 8'h00; ram[16'h19fc] = 8'h48; ram[16'h19fd] = 8'ha9; ram[16'h19fe] = 8'haa; ram[16'h19ff] = 8'h28; 

ram[16'h1a00] = 8'h9c; ram[16'h1a01] = 8'h05; ram[16'h1a02] = 8'h02; ram[16'h1a03] = 8'h9c; ram[16'h1a04] = 8'h06; ram[16'h1a05] = 8'h02; ram[16'h1a06] = 8'h9c; ram[16'h1a07] = 8'h07; 
ram[16'h1a08] = 8'h02; ram[16'h1a09] = 8'h9c; ram[16'h1a0a] = 8'h08; ram[16'h1a0b] = 8'h02; ram[16'h1a0c] = 8'h9c; ram[16'h1a0d] = 8'h09; ram[16'h1a0e] = 8'h02; ram[16'h1a0f] = 8'h08; 
ram[16'h1a10] = 8'hc9; ram[16'h1a11] = 8'haa; ram[16'h1a12] = 8'hd0; ram[16'h1a13] = 8'hfe; ram[16'h1a14] = 8'h68; ram[16'h1a15] = 8'h48; ram[16'h1a16] = 8'hc9; ram[16'h1a17] = 8'h30; 
ram[16'h1a18] = 8'hd0; ram[16'h1a19] = 8'hfe; ram[16'h1a1a] = 8'h28; ram[16'h1a1b] = 8'hbd; ram[16'h1a1c] = 8'h05; ram[16'h1a1d] = 8'h02; ram[16'h1a1e] = 8'hd0; ram[16'h1a1f] = 8'hfe; 

ram[16'h1a20] = 8'hca; ram[16'h1a21] = 8'h10; ram[16'h1a22] = 8'hf8; ram[16'h1a23] = 8'ha2; ram[16'h1a24] = 8'h04; ram[16'h1a25] = 8'ha9; ram[16'h1a26] = 8'h07; ram[16'h1a27] = 8'h95; 
ram[16'h1a28] = 8'h0c; ram[16'h1a29] = 8'h0a; ram[16'h1a2a] = 8'hca; ram[16'h1a2b] = 8'h10; ram[16'h1a2c] = 8'hfa; ram[16'h1a2d] = 8'ha2; ram[16'h1a2e] = 8'h04; ram[16'h1a2f] = 8'ha9; 
ram[16'h1a30] = 8'hff; ram[16'h1a31] = 8'h48; ram[16'h1a32] = 8'ha9; ram[16'h1a33] = 8'h55; ram[16'h1a34] = 8'h28; ram[16'h1a35] = 8'h74; ram[16'h1a36] = 8'h0c; ram[16'h1a37] = 8'h08; 
ram[16'h1a38] = 8'hc9; ram[16'h1a39] = 8'h55; ram[16'h1a3a] = 8'hd0; ram[16'h1a3b] = 8'hfe; ram[16'h1a3c] = 8'h68; ram[16'h1a3d] = 8'h48; ram[16'h1a3e] = 8'hc9; ram[16'h1a3f] = 8'hff; 

ram[16'h1a40] = 8'hd0; ram[16'h1a41] = 8'hfe; ram[16'h1a42] = 8'h28; ram[16'h1a43] = 8'hca; ram[16'h1a44] = 8'h10; ram[16'h1a45] = 8'he9; ram[16'h1a46] = 8'ha2; ram[16'h1a47] = 8'h04; 
ram[16'h1a48] = 8'hb5; ram[16'h1a49] = 8'h0c; ram[16'h1a4a] = 8'hd0; ram[16'h1a4b] = 8'hfe; ram[16'h1a4c] = 8'hca; ram[16'h1a4d] = 8'h10; ram[16'h1a4e] = 8'hf9; ram[16'h1a4f] = 8'ha2; 
ram[16'h1a50] = 8'h04; ram[16'h1a51] = 8'ha9; ram[16'h1a52] = 8'h07; ram[16'h1a53] = 8'h95; ram[16'h1a54] = 8'h0c; ram[16'h1a55] = 8'h0a; ram[16'h1a56] = 8'hca; ram[16'h1a57] = 8'h10; 
ram[16'h1a58] = 8'hfa; ram[16'h1a59] = 8'ha2; ram[16'h1a5a] = 8'h04; ram[16'h1a5b] = 8'ha9; ram[16'h1a5c] = 8'h00; ram[16'h1a5d] = 8'h48; ram[16'h1a5e] = 8'ha9; ram[16'h1a5f] = 8'haa; 

ram[16'h1a60] = 8'h28; ram[16'h1a61] = 8'h74; ram[16'h1a62] = 8'h0c; ram[16'h1a63] = 8'h08; ram[16'h1a64] = 8'hc9; ram[16'h1a65] = 8'haa; ram[16'h1a66] = 8'hd0; ram[16'h1a67] = 8'hfe; 
ram[16'h1a68] = 8'h68; ram[16'h1a69] = 8'h48; ram[16'h1a6a] = 8'hc9; ram[16'h1a6b] = 8'h30; ram[16'h1a6c] = 8'hd0; ram[16'h1a6d] = 8'hfe; ram[16'h1a6e] = 8'h28; ram[16'h1a6f] = 8'hca; 
ram[16'h1a70] = 8'h10; ram[16'h1a71] = 8'he9; ram[16'h1a72] = 8'ha2; ram[16'h1a73] = 8'h04; ram[16'h1a74] = 8'hb5; ram[16'h1a75] = 8'h0c; ram[16'h1a76] = 8'hd0; ram[16'h1a77] = 8'hfe; 
ram[16'h1a78] = 8'hca; ram[16'h1a79] = 8'h10; ram[16'h1a7a] = 8'hf9; ram[16'h1a7b] = 8'ha2; ram[16'h1a7c] = 8'h04; ram[16'h1a7d] = 8'ha9; ram[16'h1a7e] = 8'h07; ram[16'h1a7f] = 8'h9d; 

ram[16'h1a80] = 8'h05; ram[16'h1a81] = 8'h02; ram[16'h1a82] = 8'h0a; ram[16'h1a83] = 8'hca; ram[16'h1a84] = 8'h10; ram[16'h1a85] = 8'hf9; ram[16'h1a86] = 8'ha2; ram[16'h1a87] = 8'h04; 
ram[16'h1a88] = 8'ha9; ram[16'h1a89] = 8'hff; ram[16'h1a8a] = 8'h48; ram[16'h1a8b] = 8'ha9; ram[16'h1a8c] = 8'h55; ram[16'h1a8d] = 8'h28; ram[16'h1a8e] = 8'h9e; ram[16'h1a8f] = 8'h05; 
ram[16'h1a90] = 8'h02; ram[16'h1a91] = 8'h08; ram[16'h1a92] = 8'hc9; ram[16'h1a93] = 8'h55; ram[16'h1a94] = 8'hd0; ram[16'h1a95] = 8'hfe; ram[16'h1a96] = 8'h68; ram[16'h1a97] = 8'h48; 
ram[16'h1a98] = 8'hc9; ram[16'h1a99] = 8'hff; ram[16'h1a9a] = 8'hd0; ram[16'h1a9b] = 8'hfe; ram[16'h1a9c] = 8'h28; ram[16'h1a9d] = 8'hca; ram[16'h1a9e] = 8'h10; ram[16'h1a9f] = 8'he8; 

ram[16'h1aa0] = 8'ha2; ram[16'h1aa1] = 8'h04; ram[16'h1aa2] = 8'hbd; ram[16'h1aa3] = 8'h05; ram[16'h1aa4] = 8'h02; ram[16'h1aa5] = 8'hd0; ram[16'h1aa6] = 8'hfe; ram[16'h1aa7] = 8'hca; 
ram[16'h1aa8] = 8'h10; ram[16'h1aa9] = 8'hf8; ram[16'h1aaa] = 8'ha2; ram[16'h1aab] = 8'h04; ram[16'h1aac] = 8'ha9; ram[16'h1aad] = 8'h07; ram[16'h1aae] = 8'h9d; ram[16'h1aaf] = 8'h05; 
ram[16'h1ab0] = 8'h02; ram[16'h1ab1] = 8'h0a; ram[16'h1ab2] = 8'hca; ram[16'h1ab3] = 8'h10; ram[16'h1ab4] = 8'hf9; ram[16'h1ab5] = 8'ha2; ram[16'h1ab6] = 8'h04; ram[16'h1ab7] = 8'ha9; 
ram[16'h1ab8] = 8'h00; ram[16'h1ab9] = 8'h48; ram[16'h1aba] = 8'ha9; ram[16'h1abb] = 8'haa; ram[16'h1abc] = 8'h28; ram[16'h1abd] = 8'h9e; ram[16'h1abe] = 8'h05; ram[16'h1abf] = 8'h02; 

ram[16'h1ac0] = 8'h08; ram[16'h1ac1] = 8'hc9; ram[16'h1ac2] = 8'haa; ram[16'h1ac3] = 8'hd0; ram[16'h1ac4] = 8'hfe; ram[16'h1ac5] = 8'h68; ram[16'h1ac6] = 8'h48; ram[16'h1ac7] = 8'hc9; 
ram[16'h1ac8] = 8'h30; ram[16'h1ac9] = 8'hd0; ram[16'h1aca] = 8'hfe; ram[16'h1acb] = 8'h28; ram[16'h1acc] = 8'hca; ram[16'h1acd] = 8'h10; ram[16'h1ace] = 8'he8; ram[16'h1acf] = 8'ha2; 
ram[16'h1ad0] = 8'h04; ram[16'h1ad1] = 8'hbd; ram[16'h1ad2] = 8'h05; ram[16'h1ad3] = 8'h02; ram[16'h1ad4] = 8'hd0; ram[16'h1ad5] = 8'hfe; ram[16'h1ad6] = 8'hca; ram[16'h1ad7] = 8'h10; 
ram[16'h1ad8] = 8'hf8; ram[16'h1ad9] = 8'hc0; ram[16'h1ada] = 8'h7b; ram[16'h1adb] = 8'hd0; ram[16'h1adc] = 8'hfe; ram[16'h1add] = 8'hba; ram[16'h1ade] = 8'he0; ram[16'h1adf] = 8'hff; 

ram[16'h1ae0] = 8'hd0; ram[16'h1ae1] = 8'hfe; ram[16'h1ae2] = 8'had; ram[16'h1ae3] = 8'h02; ram[16'h1ae4] = 8'h02; ram[16'h1ae5] = 8'hc9; ram[16'h1ae6] = 8'h0e; ram[16'h1ae7] = 8'hd0; 
ram[16'h1ae8] = 8'hfe; ram[16'h1ae9] = 8'ha9; ram[16'h1aea] = 8'h0f; ram[16'h1aeb] = 8'h8d; ram[16'h1aec] = 8'h02; ram[16'h1aed] = 8'h02; ram[16'h1aee] = 8'ha0; ram[16'h1aef] = 8'h42; 
ram[16'h1af0] = 8'ha2; ram[16'h1af1] = 8'h03; ram[16'h1af2] = 8'ha9; ram[16'h1af3] = 8'h00; ram[16'h1af4] = 8'h48; ram[16'h1af5] = 8'ha9; ram[16'h1af6] = 8'hff; ram[16'h1af7] = 8'h28; 
ram[16'h1af8] = 8'h34; ram[16'h1af9] = 8'h13; ram[16'h1afa] = 8'h08; ram[16'h1afb] = 8'hc9; ram[16'h1afc] = 8'hff; ram[16'h1afd] = 8'hd0; ram[16'h1afe] = 8'hfe; ram[16'h1aff] = 8'h68; 

ram[16'h1b00] = 8'h48; ram[16'h1b01] = 8'hc9; ram[16'h1b02] = 8'h32; ram[16'h1b03] = 8'hd0; ram[16'h1b04] = 8'hfe; ram[16'h1b05] = 8'h28; ram[16'h1b06] = 8'hca; ram[16'h1b07] = 8'ha9; 
ram[16'h1b08] = 8'h00; ram[16'h1b09] = 8'h48; ram[16'h1b0a] = 8'ha9; ram[16'h1b0b] = 8'h01; ram[16'h1b0c] = 8'h28; ram[16'h1b0d] = 8'h34; ram[16'h1b0e] = 8'h13; ram[16'h1b0f] = 8'h08; 
ram[16'h1b10] = 8'hc9; ram[16'h1b11] = 8'h01; ram[16'h1b12] = 8'hd0; ram[16'h1b13] = 8'hfe; ram[16'h1b14] = 8'h68; ram[16'h1b15] = 8'h48; ram[16'h1b16] = 8'hc9; ram[16'h1b17] = 8'h70; 
ram[16'h1b18] = 8'hd0; ram[16'h1b19] = 8'hfe; ram[16'h1b1a] = 8'h28; ram[16'h1b1b] = 8'hca; ram[16'h1b1c] = 8'ha9; ram[16'h1b1d] = 8'h00; ram[16'h1b1e] = 8'h48; ram[16'h1b1f] = 8'ha9; 

ram[16'h1b20] = 8'h01; ram[16'h1b21] = 8'h28; ram[16'h1b22] = 8'h34; ram[16'h1b23] = 8'h13; ram[16'h1b24] = 8'h08; ram[16'h1b25] = 8'hc9; ram[16'h1b26] = 8'h01; ram[16'h1b27] = 8'hd0; 
ram[16'h1b28] = 8'hfe; ram[16'h1b29] = 8'h68; ram[16'h1b2a] = 8'h48; ram[16'h1b2b] = 8'hc9; ram[16'h1b2c] = 8'hb2; ram[16'h1b2d] = 8'hd0; ram[16'h1b2e] = 8'hfe; ram[16'h1b2f] = 8'h28; 
ram[16'h1b30] = 8'hca; ram[16'h1b31] = 8'ha9; ram[16'h1b32] = 8'h00; ram[16'h1b33] = 8'h48; ram[16'h1b34] = 8'ha9; ram[16'h1b35] = 8'h01; ram[16'h1b36] = 8'h28; ram[16'h1b37] = 8'h34; 
ram[16'h1b38] = 8'h13; ram[16'h1b39] = 8'h08; ram[16'h1b3a] = 8'hc9; ram[16'h1b3b] = 8'h01; ram[16'h1b3c] = 8'hd0; ram[16'h1b3d] = 8'hfe; ram[16'h1b3e] = 8'h68; ram[16'h1b3f] = 8'h48; 

ram[16'h1b40] = 8'hc9; ram[16'h1b41] = 8'hf0; ram[16'h1b42] = 8'hd0; ram[16'h1b43] = 8'hfe; ram[16'h1b44] = 8'h28; ram[16'h1b45] = 8'ha9; ram[16'h1b46] = 8'hff; ram[16'h1b47] = 8'h48; 
ram[16'h1b48] = 8'ha9; ram[16'h1b49] = 8'h01; ram[16'h1b4a] = 8'h28; ram[16'h1b4b] = 8'h34; ram[16'h1b4c] = 8'h13; ram[16'h1b4d] = 8'h08; ram[16'h1b4e] = 8'hc9; ram[16'h1b4f] = 8'h01; 
ram[16'h1b50] = 8'hd0; ram[16'h1b51] = 8'hfe; ram[16'h1b52] = 8'h68; ram[16'h1b53] = 8'h48; ram[16'h1b54] = 8'hc9; ram[16'h1b55] = 8'hfd; ram[16'h1b56] = 8'hd0; ram[16'h1b57] = 8'hfe; 
ram[16'h1b58] = 8'h28; ram[16'h1b59] = 8'he8; ram[16'h1b5a] = 8'ha9; ram[16'h1b5b] = 8'hff; ram[16'h1b5c] = 8'h48; ram[16'h1b5d] = 8'ha9; ram[16'h1b5e] = 8'h01; ram[16'h1b5f] = 8'h28; 

ram[16'h1b60] = 8'h34; ram[16'h1b61] = 8'h13; ram[16'h1b62] = 8'h08; ram[16'h1b63] = 8'hc9; ram[16'h1b64] = 8'h01; ram[16'h1b65] = 8'hd0; ram[16'h1b66] = 8'hfe; ram[16'h1b67] = 8'h68; 
ram[16'h1b68] = 8'h48; ram[16'h1b69] = 8'hc9; ram[16'h1b6a] = 8'hbf; ram[16'h1b6b] = 8'hd0; ram[16'h1b6c] = 8'hfe; ram[16'h1b6d] = 8'h28; ram[16'h1b6e] = 8'he8; ram[16'h1b6f] = 8'ha9; 
ram[16'h1b70] = 8'hff; ram[16'h1b71] = 8'h48; ram[16'h1b72] = 8'ha9; ram[16'h1b73] = 8'h01; ram[16'h1b74] = 8'h28; ram[16'h1b75] = 8'h34; ram[16'h1b76] = 8'h13; ram[16'h1b77] = 8'h08; 
ram[16'h1b78] = 8'hc9; ram[16'h1b79] = 8'h01; ram[16'h1b7a] = 8'hd0; ram[16'h1b7b] = 8'hfe; ram[16'h1b7c] = 8'h68; ram[16'h1b7d] = 8'h48; ram[16'h1b7e] = 8'hc9; ram[16'h1b7f] = 8'h7d; 

ram[16'h1b80] = 8'hd0; ram[16'h1b81] = 8'hfe; ram[16'h1b82] = 8'h28; ram[16'h1b83] = 8'he8; ram[16'h1b84] = 8'ha9; ram[16'h1b85] = 8'hff; ram[16'h1b86] = 8'h48; ram[16'h1b87] = 8'ha9; 
ram[16'h1b88] = 8'hff; ram[16'h1b89] = 8'h28; ram[16'h1b8a] = 8'h34; ram[16'h1b8b] = 8'h13; ram[16'h1b8c] = 8'h08; ram[16'h1b8d] = 8'hc9; ram[16'h1b8e] = 8'hff; ram[16'h1b8f] = 8'hd0; 
ram[16'h1b90] = 8'hfe; ram[16'h1b91] = 8'h68; ram[16'h1b92] = 8'h48; ram[16'h1b93] = 8'hc9; ram[16'h1b94] = 8'h3f; ram[16'h1b95] = 8'hd0; ram[16'h1b96] = 8'hfe; ram[16'h1b97] = 8'h28; 
ram[16'h1b98] = 8'ha9; ram[16'h1b99] = 8'h00; ram[16'h1b9a] = 8'h48; ram[16'h1b9b] = 8'ha9; ram[16'h1b9c] = 8'hff; ram[16'h1b9d] = 8'h28; ram[16'h1b9e] = 8'h3c; ram[16'h1b9f] = 8'h10; 

ram[16'h1ba0] = 8'h02; ram[16'h1ba1] = 8'h08; ram[16'h1ba2] = 8'hc9; ram[16'h1ba3] = 8'hff; ram[16'h1ba4] = 8'hd0; ram[16'h1ba5] = 8'hfe; ram[16'h1ba6] = 8'h68; ram[16'h1ba7] = 8'h48; 
ram[16'h1ba8] = 8'hc9; ram[16'h1ba9] = 8'h32; ram[16'h1baa] = 8'hd0; ram[16'h1bab] = 8'hfe; ram[16'h1bac] = 8'h28; ram[16'h1bad] = 8'hca; ram[16'h1bae] = 8'ha9; ram[16'h1baf] = 8'h00; 
ram[16'h1bb0] = 8'h48; ram[16'h1bb1] = 8'ha9; ram[16'h1bb2] = 8'h01; ram[16'h1bb3] = 8'h28; ram[16'h1bb4] = 8'h3c; ram[16'h1bb5] = 8'h10; ram[16'h1bb6] = 8'h02; ram[16'h1bb7] = 8'h08; 
ram[16'h1bb8] = 8'hc9; ram[16'h1bb9] = 8'h01; ram[16'h1bba] = 8'hd0; ram[16'h1bbb] = 8'hfe; ram[16'h1bbc] = 8'h68; ram[16'h1bbd] = 8'h48; ram[16'h1bbe] = 8'hc9; ram[16'h1bbf] = 8'h70; 

ram[16'h1bc0] = 8'hd0; ram[16'h1bc1] = 8'hfe; ram[16'h1bc2] = 8'h28; ram[16'h1bc3] = 8'hca; ram[16'h1bc4] = 8'ha9; ram[16'h1bc5] = 8'h00; ram[16'h1bc6] = 8'h48; ram[16'h1bc7] = 8'ha9; 
ram[16'h1bc8] = 8'h01; ram[16'h1bc9] = 8'h28; ram[16'h1bca] = 8'h3c; ram[16'h1bcb] = 8'h10; ram[16'h1bcc] = 8'h02; ram[16'h1bcd] = 8'h08; ram[16'h1bce] = 8'hc9; ram[16'h1bcf] = 8'h01; 
ram[16'h1bd0] = 8'hd0; ram[16'h1bd1] = 8'hfe; ram[16'h1bd2] = 8'h68; ram[16'h1bd3] = 8'h48; ram[16'h1bd4] = 8'hc9; ram[16'h1bd5] = 8'hb2; ram[16'h1bd6] = 8'hd0; ram[16'h1bd7] = 8'hfe; 
ram[16'h1bd8] = 8'h28; ram[16'h1bd9] = 8'hca; ram[16'h1bda] = 8'ha9; ram[16'h1bdb] = 8'h00; ram[16'h1bdc] = 8'h48; ram[16'h1bdd] = 8'ha9; ram[16'h1bde] = 8'h01; ram[16'h1bdf] = 8'h28; 

ram[16'h1be0] = 8'h3c; ram[16'h1be1] = 8'h10; ram[16'h1be2] = 8'h02; ram[16'h1be3] = 8'h08; ram[16'h1be4] = 8'hc9; ram[16'h1be5] = 8'h01; ram[16'h1be6] = 8'hd0; ram[16'h1be7] = 8'hfe; 
ram[16'h1be8] = 8'h68; ram[16'h1be9] = 8'h48; ram[16'h1bea] = 8'hc9; ram[16'h1beb] = 8'hf0; ram[16'h1bec] = 8'hd0; ram[16'h1bed] = 8'hfe; ram[16'h1bee] = 8'h28; ram[16'h1bef] = 8'ha9; 
ram[16'h1bf0] = 8'hff; ram[16'h1bf1] = 8'h48; ram[16'h1bf2] = 8'ha9; ram[16'h1bf3] = 8'h01; ram[16'h1bf4] = 8'h28; ram[16'h1bf5] = 8'h3c; ram[16'h1bf6] = 8'h10; ram[16'h1bf7] = 8'h02; 
ram[16'h1bf8] = 8'h08; ram[16'h1bf9] = 8'hc9; ram[16'h1bfa] = 8'h01; ram[16'h1bfb] = 8'hd0; ram[16'h1bfc] = 8'hfe; ram[16'h1bfd] = 8'h68; ram[16'h1bfe] = 8'h48; ram[16'h1bff] = 8'hc9; 

ram[16'h1c00] = 8'hfd; ram[16'h1c01] = 8'hd0; ram[16'h1c02] = 8'hfe; ram[16'h1c03] = 8'h28; ram[16'h1c04] = 8'he8; ram[16'h1c05] = 8'ha9; ram[16'h1c06] = 8'hff; ram[16'h1c07] = 8'h48; 
ram[16'h1c08] = 8'ha9; ram[16'h1c09] = 8'h01; ram[16'h1c0a] = 8'h28; ram[16'h1c0b] = 8'h3c; ram[16'h1c0c] = 8'h10; ram[16'h1c0d] = 8'h02; ram[16'h1c0e] = 8'h08; ram[16'h1c0f] = 8'hc9; 
ram[16'h1c10] = 8'h01; ram[16'h1c11] = 8'hd0; ram[16'h1c12] = 8'hfe; ram[16'h1c13] = 8'h68; ram[16'h1c14] = 8'h48; ram[16'h1c15] = 8'hc9; ram[16'h1c16] = 8'hbf; ram[16'h1c17] = 8'hd0; 
ram[16'h1c18] = 8'hfe; ram[16'h1c19] = 8'h28; ram[16'h1c1a] = 8'he8; ram[16'h1c1b] = 8'ha9; ram[16'h1c1c] = 8'hff; ram[16'h1c1d] = 8'h48; ram[16'h1c1e] = 8'ha9; ram[16'h1c1f] = 8'h01; 

ram[16'h1c20] = 8'h28; ram[16'h1c21] = 8'h3c; ram[16'h1c22] = 8'h10; ram[16'h1c23] = 8'h02; ram[16'h1c24] = 8'h08; ram[16'h1c25] = 8'hc9; ram[16'h1c26] = 8'h01; ram[16'h1c27] = 8'hd0; 
ram[16'h1c28] = 8'hfe; ram[16'h1c29] = 8'h68; ram[16'h1c2a] = 8'h48; ram[16'h1c2b] = 8'hc9; ram[16'h1c2c] = 8'h7d; ram[16'h1c2d] = 8'hd0; ram[16'h1c2e] = 8'hfe; ram[16'h1c2f] = 8'h28; 
ram[16'h1c30] = 8'he8; ram[16'h1c31] = 8'ha9; ram[16'h1c32] = 8'hff; ram[16'h1c33] = 8'h48; ram[16'h1c34] = 8'ha9; ram[16'h1c35] = 8'hff; ram[16'h1c36] = 8'h28; ram[16'h1c37] = 8'h3c; 
ram[16'h1c38] = 8'h10; ram[16'h1c39] = 8'h02; ram[16'h1c3a] = 8'h08; ram[16'h1c3b] = 8'hc9; ram[16'h1c3c] = 8'hff; ram[16'h1c3d] = 8'hd0; ram[16'h1c3e] = 8'hfe; ram[16'h1c3f] = 8'h68; 

ram[16'h1c40] = 8'h48; ram[16'h1c41] = 8'hc9; ram[16'h1c42] = 8'h3f; ram[16'h1c43] = 8'hd0; ram[16'h1c44] = 8'hfe; ram[16'h1c45] = 8'h28; ram[16'h1c46] = 8'ha9; ram[16'h1c47] = 8'h00; 
ram[16'h1c48] = 8'h48; ram[16'h1c49] = 8'ha9; ram[16'h1c4a] = 8'hff; ram[16'h1c4b] = 8'h28; ram[16'h1c4c] = 8'h89; ram[16'h1c4d] = 8'h00; ram[16'h1c4e] = 8'h08; ram[16'h1c4f] = 8'hc9; 
ram[16'h1c50] = 8'hff; ram[16'h1c51] = 8'hd0; ram[16'h1c52] = 8'hfe; ram[16'h1c53] = 8'h68; ram[16'h1c54] = 8'h48; ram[16'h1c55] = 8'hc9; ram[16'h1c56] = 8'h32; ram[16'h1c57] = 8'hd0; 
ram[16'h1c58] = 8'hfe; ram[16'h1c59] = 8'h28; ram[16'h1c5a] = 8'hca; ram[16'h1c5b] = 8'ha9; ram[16'h1c5c] = 8'h00; ram[16'h1c5d] = 8'h48; ram[16'h1c5e] = 8'ha9; ram[16'h1c5f] = 8'h01; 

ram[16'h1c60] = 8'h28; ram[16'h1c61] = 8'h89; ram[16'h1c62] = 8'h41; ram[16'h1c63] = 8'h08; ram[16'h1c64] = 8'hc9; ram[16'h1c65] = 8'h01; ram[16'h1c66] = 8'hd0; ram[16'h1c67] = 8'hfe; 
ram[16'h1c68] = 8'h68; ram[16'h1c69] = 8'h48; ram[16'h1c6a] = 8'hc9; ram[16'h1c6b] = 8'h30; ram[16'h1c6c] = 8'hd0; ram[16'h1c6d] = 8'hfe; ram[16'h1c6e] = 8'h28; ram[16'h1c6f] = 8'hca; 
ram[16'h1c70] = 8'ha9; ram[16'h1c71] = 8'h00; ram[16'h1c72] = 8'h48; ram[16'h1c73] = 8'ha9; ram[16'h1c74] = 8'h01; ram[16'h1c75] = 8'h28; ram[16'h1c76] = 8'h89; ram[16'h1c77] = 8'h82; 
ram[16'h1c78] = 8'h08; ram[16'h1c79] = 8'hc9; ram[16'h1c7a] = 8'h01; ram[16'h1c7b] = 8'hd0; ram[16'h1c7c] = 8'hfe; ram[16'h1c7d] = 8'h68; ram[16'h1c7e] = 8'h48; ram[16'h1c7f] = 8'hc9; 

ram[16'h1c80] = 8'h32; ram[16'h1c81] = 8'hd0; ram[16'h1c82] = 8'hfe; ram[16'h1c83] = 8'h28; ram[16'h1c84] = 8'hca; ram[16'h1c85] = 8'ha9; ram[16'h1c86] = 8'h00; ram[16'h1c87] = 8'h48; 
ram[16'h1c88] = 8'ha9; ram[16'h1c89] = 8'h01; ram[16'h1c8a] = 8'h28; ram[16'h1c8b] = 8'h89; ram[16'h1c8c] = 8'hc3; ram[16'h1c8d] = 8'h08; ram[16'h1c8e] = 8'hc9; ram[16'h1c8f] = 8'h01; 
ram[16'h1c90] = 8'hd0; ram[16'h1c91] = 8'hfe; ram[16'h1c92] = 8'h68; ram[16'h1c93] = 8'h48; ram[16'h1c94] = 8'hc9; ram[16'h1c95] = 8'h30; ram[16'h1c96] = 8'hd0; ram[16'h1c97] = 8'hfe; 
ram[16'h1c98] = 8'h28; ram[16'h1c99] = 8'ha9; ram[16'h1c9a] = 8'hff; ram[16'h1c9b] = 8'h48; ram[16'h1c9c] = 8'ha9; ram[16'h1c9d] = 8'h01; ram[16'h1c9e] = 8'h28; ram[16'h1c9f] = 8'h89; 

ram[16'h1ca0] = 8'hc3; ram[16'h1ca1] = 8'h08; ram[16'h1ca2] = 8'hc9; ram[16'h1ca3] = 8'h01; ram[16'h1ca4] = 8'hd0; ram[16'h1ca5] = 8'hfe; ram[16'h1ca6] = 8'h68; ram[16'h1ca7] = 8'h48; 
ram[16'h1ca8] = 8'hc9; ram[16'h1ca9] = 8'hfd; ram[16'h1caa] = 8'hd0; ram[16'h1cab] = 8'hfe; ram[16'h1cac] = 8'h28; ram[16'h1cad] = 8'he8; ram[16'h1cae] = 8'ha9; ram[16'h1caf] = 8'hff; 
ram[16'h1cb0] = 8'h48; ram[16'h1cb1] = 8'ha9; ram[16'h1cb2] = 8'h01; ram[16'h1cb3] = 8'h28; ram[16'h1cb4] = 8'h89; ram[16'h1cb5] = 8'h82; ram[16'h1cb6] = 8'h08; ram[16'h1cb7] = 8'hc9; 
ram[16'h1cb8] = 8'h01; ram[16'h1cb9] = 8'hd0; ram[16'h1cba] = 8'hfe; ram[16'h1cbb] = 8'h68; ram[16'h1cbc] = 8'h48; ram[16'h1cbd] = 8'hc9; ram[16'h1cbe] = 8'hff; ram[16'h1cbf] = 8'hd0; 

ram[16'h1cc0] = 8'hfe; ram[16'h1cc1] = 8'h28; ram[16'h1cc2] = 8'he8; ram[16'h1cc3] = 8'ha9; ram[16'h1cc4] = 8'hff; ram[16'h1cc5] = 8'h48; ram[16'h1cc6] = 8'ha9; ram[16'h1cc7] = 8'h01; 
ram[16'h1cc8] = 8'h28; ram[16'h1cc9] = 8'h89; ram[16'h1cca] = 8'h41; ram[16'h1ccb] = 8'h08; ram[16'h1ccc] = 8'hc9; ram[16'h1ccd] = 8'h01; ram[16'h1cce] = 8'hd0; ram[16'h1ccf] = 8'hfe; 
ram[16'h1cd0] = 8'h68; ram[16'h1cd1] = 8'h48; ram[16'h1cd2] = 8'hc9; ram[16'h1cd3] = 8'hfd; ram[16'h1cd4] = 8'hd0; ram[16'h1cd5] = 8'hfe; ram[16'h1cd6] = 8'h28; ram[16'h1cd7] = 8'he8; 
ram[16'h1cd8] = 8'ha9; ram[16'h1cd9] = 8'hff; ram[16'h1cda] = 8'h48; ram[16'h1cdb] = 8'ha9; ram[16'h1cdc] = 8'hff; ram[16'h1cdd] = 8'h28; ram[16'h1cde] = 8'h89; ram[16'h1cdf] = 8'h00; 

ram[16'h1ce0] = 8'h08; ram[16'h1ce1] = 8'hc9; ram[16'h1ce2] = 8'hff; ram[16'h1ce3] = 8'hd0; ram[16'h1ce4] = 8'hfe; ram[16'h1ce5] = 8'h68; ram[16'h1ce6] = 8'h48; ram[16'h1ce7] = 8'hc9; 
ram[16'h1ce8] = 8'hff; ram[16'h1ce9] = 8'hd0; ram[16'h1cea] = 8'hfe; ram[16'h1ceb] = 8'h28; ram[16'h1cec] = 8'he0; ram[16'h1ced] = 8'h03; ram[16'h1cee] = 8'hd0; ram[16'h1cef] = 8'hfe; 
ram[16'h1cf0] = 8'hc0; ram[16'h1cf1] = 8'h42; ram[16'h1cf2] = 8'hd0; ram[16'h1cf3] = 8'hfe; ram[16'h1cf4] = 8'hba; ram[16'h1cf5] = 8'he0; ram[16'h1cf6] = 8'hff; ram[16'h1cf7] = 8'hd0; 
ram[16'h1cf8] = 8'hfe; ram[16'h1cf9] = 8'had; ram[16'h1cfa] = 8'h02; ram[16'h1cfb] = 8'h02; ram[16'h1cfc] = 8'hc9; ram[16'h1cfd] = 8'h0f; ram[16'h1cfe] = 8'hd0; ram[16'h1cff] = 8'hfe; 

ram[16'h1d00] = 8'ha9; ram[16'h1d01] = 8'h10; ram[16'h1d02] = 8'h8d; ram[16'h1d03] = 8'h02; ram[16'h1d04] = 8'h02; ram[16'h1d05] = 8'ha2; ram[16'h1d06] = 8'hc0; ram[16'h1d07] = 8'ha0; 
ram[16'h1d08] = 8'h00; ram[16'h1d09] = 8'h64; ram[16'h1d0a] = 8'h0d; ram[16'h1d0b] = 8'h98; ram[16'h1d0c] = 8'h25; ram[16'h1d0d] = 8'h0d; ram[16'h1d0e] = 8'h08; ram[16'h1d0f] = 8'h68; 
ram[16'h1d10] = 8'h29; ram[16'h1d11] = 8'h02; ram[16'h1d12] = 8'h85; ram[16'h1d13] = 8'h0e; ram[16'h1d14] = 8'h98; ram[16'h1d15] = 8'h49; ram[16'h1d16] = 8'hff; ram[16'h1d17] = 8'h05; 
ram[16'h1d18] = 8'h0d; ram[16'h1d19] = 8'h49; ram[16'h1d1a] = 8'hff; ram[16'h1d1b] = 8'h85; ram[16'h1d1c] = 8'h0f; ram[16'h1d1d] = 8'h98; ram[16'h1d1e] = 8'h05; ram[16'h1d1f] = 8'h0d; 

ram[16'h1d20] = 8'h85; ram[16'h1d21] = 8'h10; ram[16'h1d22] = 8'h84; ram[16'h1d23] = 8'h0c; ram[16'h1d24] = 8'ha9; ram[16'h1d25] = 8'hff; ram[16'h1d26] = 8'h48; ram[16'h1d27] = 8'ha5; 
ram[16'h1d28] = 8'h0d; ram[16'h1d29] = 8'h28; ram[16'h1d2a] = 8'h14; ram[16'h1d2b] = 8'h0c; ram[16'h1d2c] = 8'h08; ram[16'h1d2d] = 8'hc5; ram[16'h1d2e] = 8'h0d; ram[16'h1d2f] = 8'hd0; 
ram[16'h1d30] = 8'hfe; ram[16'h1d31] = 8'h68; ram[16'h1d32] = 8'h48; ram[16'h1d33] = 8'h09; ram[16'h1d34] = 8'h02; ram[16'h1d35] = 8'hc9; ram[16'h1d36] = 8'hff; ram[16'h1d37] = 8'hd0; 
ram[16'h1d38] = 8'hfe; ram[16'h1d39] = 8'h68; ram[16'h1d3a] = 8'h29; ram[16'h1d3b] = 8'h02; ram[16'h1d3c] = 8'hc5; ram[16'h1d3d] = 8'h0e; ram[16'h1d3e] = 8'hd0; ram[16'h1d3f] = 8'hfe; 

ram[16'h1d40] = 8'ha5; ram[16'h1d41] = 8'h0f; ram[16'h1d42] = 8'hc5; ram[16'h1d43] = 8'h0c; ram[16'h1d44] = 8'hd0; ram[16'h1d45] = 8'hfe; ram[16'h1d46] = 8'h8c; ram[16'h1d47] = 8'h05; 
ram[16'h1d48] = 8'h02; ram[16'h1d49] = 8'ha9; ram[16'h1d4a] = 8'hff; ram[16'h1d4b] = 8'h48; ram[16'h1d4c] = 8'ha5; ram[16'h1d4d] = 8'h0d; ram[16'h1d4e] = 8'h28; ram[16'h1d4f] = 8'h1c; 
ram[16'h1d50] = 8'h05; ram[16'h1d51] = 8'h02; ram[16'h1d52] = 8'h08; ram[16'h1d53] = 8'hc5; ram[16'h1d54] = 8'h0d; ram[16'h1d55] = 8'hd0; ram[16'h1d56] = 8'hfe; ram[16'h1d57] = 8'h68; 
ram[16'h1d58] = 8'h48; ram[16'h1d59] = 8'h09; ram[16'h1d5a] = 8'h02; ram[16'h1d5b] = 8'hc9; ram[16'h1d5c] = 8'hff; ram[16'h1d5d] = 8'hd0; ram[16'h1d5e] = 8'hfe; ram[16'h1d5f] = 8'h68; 

ram[16'h1d60] = 8'h29; ram[16'h1d61] = 8'h02; ram[16'h1d62] = 8'hc5; ram[16'h1d63] = 8'h0e; ram[16'h1d64] = 8'hd0; ram[16'h1d65] = 8'hfe; ram[16'h1d66] = 8'ha5; ram[16'h1d67] = 8'h0f; 
ram[16'h1d68] = 8'hc5; ram[16'h1d69] = 8'h0c; ram[16'h1d6a] = 8'hd0; ram[16'h1d6b] = 8'hfe; ram[16'h1d6c] = 8'h84; ram[16'h1d6d] = 8'h0c; ram[16'h1d6e] = 8'ha9; ram[16'h1d6f] = 8'h00; 
ram[16'h1d70] = 8'h48; ram[16'h1d71] = 8'ha5; ram[16'h1d72] = 8'h0d; ram[16'h1d73] = 8'h28; ram[16'h1d74] = 8'h14; ram[16'h1d75] = 8'h0c; ram[16'h1d76] = 8'h08; ram[16'h1d77] = 8'hc5; 
ram[16'h1d78] = 8'h0d; ram[16'h1d79] = 8'hd0; ram[16'h1d7a] = 8'hfe; ram[16'h1d7b] = 8'h68; ram[16'h1d7c] = 8'h48; ram[16'h1d7d] = 8'h09; ram[16'h1d7e] = 8'h02; ram[16'h1d7f] = 8'hc9; 

ram[16'h1d80] = 8'h32; ram[16'h1d81] = 8'hd0; ram[16'h1d82] = 8'hfe; ram[16'h1d83] = 8'h68; ram[16'h1d84] = 8'h29; ram[16'h1d85] = 8'h02; ram[16'h1d86] = 8'hc5; ram[16'h1d87] = 8'h0e; 
ram[16'h1d88] = 8'hd0; ram[16'h1d89] = 8'hfe; ram[16'h1d8a] = 8'ha5; ram[16'h1d8b] = 8'h0f; ram[16'h1d8c] = 8'hc5; ram[16'h1d8d] = 8'h0c; ram[16'h1d8e] = 8'hd0; ram[16'h1d8f] = 8'hfe; 
ram[16'h1d90] = 8'h8c; ram[16'h1d91] = 8'h05; ram[16'h1d92] = 8'h02; ram[16'h1d93] = 8'ha9; ram[16'h1d94] = 8'h00; ram[16'h1d95] = 8'h48; ram[16'h1d96] = 8'ha5; ram[16'h1d97] = 8'h0d; 
ram[16'h1d98] = 8'h28; ram[16'h1d99] = 8'h1c; ram[16'h1d9a] = 8'h05; ram[16'h1d9b] = 8'h02; ram[16'h1d9c] = 8'h08; ram[16'h1d9d] = 8'hc5; ram[16'h1d9e] = 8'h0d; ram[16'h1d9f] = 8'hd0; 

ram[16'h1da0] = 8'hfe; ram[16'h1da1] = 8'h68; ram[16'h1da2] = 8'h48; ram[16'h1da3] = 8'h09; ram[16'h1da4] = 8'h02; ram[16'h1da5] = 8'hc9; ram[16'h1da6] = 8'h32; ram[16'h1da7] = 8'hd0; 
ram[16'h1da8] = 8'hfe; ram[16'h1da9] = 8'h68; ram[16'h1daa] = 8'h29; ram[16'h1dab] = 8'h02; ram[16'h1dac] = 8'hc5; ram[16'h1dad] = 8'h0e; ram[16'h1dae] = 8'hd0; ram[16'h1daf] = 8'hfe; 
ram[16'h1db0] = 8'ha5; ram[16'h1db1] = 8'h0f; ram[16'h1db2] = 8'hc5; ram[16'h1db3] = 8'h0c; ram[16'h1db4] = 8'hd0; ram[16'h1db5] = 8'hfe; ram[16'h1db6] = 8'h84; ram[16'h1db7] = 8'h0c; 
ram[16'h1db8] = 8'ha9; ram[16'h1db9] = 8'hff; ram[16'h1dba] = 8'h48; ram[16'h1dbb] = 8'ha5; ram[16'h1dbc] = 8'h0d; ram[16'h1dbd] = 8'h28; ram[16'h1dbe] = 8'h04; ram[16'h1dbf] = 8'h0c; 

ram[16'h1dc0] = 8'h08; ram[16'h1dc1] = 8'hc5; ram[16'h1dc2] = 8'h0d; ram[16'h1dc3] = 8'hd0; ram[16'h1dc4] = 8'hfe; ram[16'h1dc5] = 8'h68; ram[16'h1dc6] = 8'h48; ram[16'h1dc7] = 8'h09; 
ram[16'h1dc8] = 8'h02; ram[16'h1dc9] = 8'hc9; ram[16'h1dca] = 8'hff; ram[16'h1dcb] = 8'hd0; ram[16'h1dcc] = 8'hfe; ram[16'h1dcd] = 8'h68; ram[16'h1dce] = 8'h29; ram[16'h1dcf] = 8'h02; 
ram[16'h1dd0] = 8'hc5; ram[16'h1dd1] = 8'h0e; ram[16'h1dd2] = 8'hd0; ram[16'h1dd3] = 8'hfe; ram[16'h1dd4] = 8'ha5; ram[16'h1dd5] = 8'h10; ram[16'h1dd6] = 8'hc5; ram[16'h1dd7] = 8'h0c; 
ram[16'h1dd8] = 8'hd0; ram[16'h1dd9] = 8'hfe; ram[16'h1dda] = 8'h8c; ram[16'h1ddb] = 8'h05; ram[16'h1ddc] = 8'h02; ram[16'h1ddd] = 8'ha9; ram[16'h1dde] = 8'hff; ram[16'h1ddf] = 8'h48; 

ram[16'h1de0] = 8'ha5; ram[16'h1de1] = 8'h0d; ram[16'h1de2] = 8'h28; ram[16'h1de3] = 8'h0c; ram[16'h1de4] = 8'h05; ram[16'h1de5] = 8'h02; ram[16'h1de6] = 8'h08; ram[16'h1de7] = 8'hc5; 
ram[16'h1de8] = 8'h0d; ram[16'h1de9] = 8'hd0; ram[16'h1dea] = 8'hfe; ram[16'h1deb] = 8'h68; ram[16'h1dec] = 8'h48; ram[16'h1ded] = 8'h09; ram[16'h1dee] = 8'h02; ram[16'h1def] = 8'hc9; 
ram[16'h1df0] = 8'hff; ram[16'h1df1] = 8'hd0; ram[16'h1df2] = 8'hfe; ram[16'h1df3] = 8'h68; ram[16'h1df4] = 8'h29; ram[16'h1df5] = 8'h02; ram[16'h1df6] = 8'hc5; ram[16'h1df7] = 8'h0e; 
ram[16'h1df8] = 8'hd0; ram[16'h1df9] = 8'hfe; ram[16'h1dfa] = 8'ha5; ram[16'h1dfb] = 8'h10; ram[16'h1dfc] = 8'hc5; ram[16'h1dfd] = 8'h0c; ram[16'h1dfe] = 8'hd0; ram[16'h1dff] = 8'hfe; 

ram[16'h1e00] = 8'h84; ram[16'h1e01] = 8'h0c; ram[16'h1e02] = 8'ha9; ram[16'h1e03] = 8'h00; ram[16'h1e04] = 8'h48; ram[16'h1e05] = 8'ha5; ram[16'h1e06] = 8'h0d; ram[16'h1e07] = 8'h28; 
ram[16'h1e08] = 8'h04; ram[16'h1e09] = 8'h0c; ram[16'h1e0a] = 8'h08; ram[16'h1e0b] = 8'hc5; ram[16'h1e0c] = 8'h0d; ram[16'h1e0d] = 8'hd0; ram[16'h1e0e] = 8'hfe; ram[16'h1e0f] = 8'h68; 
ram[16'h1e10] = 8'h48; ram[16'h1e11] = 8'h09; ram[16'h1e12] = 8'h02; ram[16'h1e13] = 8'hc9; ram[16'h1e14] = 8'h32; ram[16'h1e15] = 8'hd0; ram[16'h1e16] = 8'hfe; ram[16'h1e17] = 8'h68; 
ram[16'h1e18] = 8'h29; ram[16'h1e19] = 8'h02; ram[16'h1e1a] = 8'hc5; ram[16'h1e1b] = 8'h0e; ram[16'h1e1c] = 8'hd0; ram[16'h1e1d] = 8'hfe; ram[16'h1e1e] = 8'ha5; ram[16'h1e1f] = 8'h10; 

ram[16'h1e20] = 8'hc5; ram[16'h1e21] = 8'h0c; ram[16'h1e22] = 8'hd0; ram[16'h1e23] = 8'hfe; ram[16'h1e24] = 8'h8c; ram[16'h1e25] = 8'h05; ram[16'h1e26] = 8'h02; ram[16'h1e27] = 8'ha9; 
ram[16'h1e28] = 8'h00; ram[16'h1e29] = 8'h48; ram[16'h1e2a] = 8'ha5; ram[16'h1e2b] = 8'h0d; ram[16'h1e2c] = 8'h28; ram[16'h1e2d] = 8'h0c; ram[16'h1e2e] = 8'h05; ram[16'h1e2f] = 8'h02; 
ram[16'h1e30] = 8'h08; ram[16'h1e31] = 8'hc5; ram[16'h1e32] = 8'h0d; ram[16'h1e33] = 8'hd0; ram[16'h1e34] = 8'hfe; ram[16'h1e35] = 8'h68; ram[16'h1e36] = 8'h48; ram[16'h1e37] = 8'h09; 
ram[16'h1e38] = 8'h02; ram[16'h1e39] = 8'hc9; ram[16'h1e3a] = 8'h32; ram[16'h1e3b] = 8'hd0; ram[16'h1e3c] = 8'hfe; ram[16'h1e3d] = 8'h68; ram[16'h1e3e] = 8'h29; ram[16'h1e3f] = 8'h02; 

ram[16'h1e40] = 8'hc5; ram[16'h1e41] = 8'h0e; ram[16'h1e42] = 8'hd0; ram[16'h1e43] = 8'hfe; ram[16'h1e44] = 8'ha5; ram[16'h1e45] = 8'h10; ram[16'h1e46] = 8'hc5; ram[16'h1e47] = 8'h0c; 
ram[16'h1e48] = 8'hd0; ram[16'h1e49] = 8'hfe; ram[16'h1e4a] = 8'hc8; ram[16'h1e4b] = 8'hd0; ram[16'h1e4c] = 8'h04; ram[16'h1e4d] = 8'he6; ram[16'h1e4e] = 8'h0d; ram[16'h1e4f] = 8'hf0; 
ram[16'h1e50] = 8'h03; ram[16'h1e51] = 8'h4c; ram[16'h1e52] = 8'h0b; ram[16'h1e53] = 8'h1d; ram[16'h1e54] = 8'he0; ram[16'h1e55] = 8'hc0; ram[16'h1e56] = 8'hd0; ram[16'h1e57] = 8'hfe; 
ram[16'h1e58] = 8'hba; ram[16'h1e59] = 8'he0; ram[16'h1e5a] = 8'hff; ram[16'h1e5b] = 8'hd0; ram[16'h1e5c] = 8'hfe; ram[16'h1e5d] = 8'had; ram[16'h1e5e] = 8'h02; ram[16'h1e5f] = 8'h02; 

ram[16'h1e60] = 8'hc9; ram[16'h1e61] = 8'h10; ram[16'h1e62] = 8'hd0; ram[16'h1e63] = 8'hfe; ram[16'h1e64] = 8'ha9; ram[16'h1e65] = 8'h11; ram[16'h1e66] = 8'h8d; ram[16'h1e67] = 8'h02; 
ram[16'h1e68] = 8'h02; ram[16'h1e69] = 8'ha2; ram[16'h1e6a] = 8'hba; ram[16'h1e6b] = 8'ha0; ram[16'h1e6c] = 8'hd0; ram[16'h1e6d] = 8'ha9; ram[16'h1e6e] = 8'hff; ram[16'h1e6f] = 8'h85; 
ram[16'h1e70] = 8'h0c; ram[16'h1e71] = 8'ha9; ram[16'h1e72] = 8'h00; ram[16'h1e73] = 8'h48; ram[16'h1e74] = 8'ha9; ram[16'h1e75] = 8'ha5; ram[16'h1e76] = 8'h28; ram[16'h1e77] = 8'h07; 
ram[16'h1e78] = 8'h0c; ram[16'h1e79] = 8'h08; ram[16'h1e7a] = 8'hc9; ram[16'h1e7b] = 8'ha5; ram[16'h1e7c] = 8'hd0; ram[16'h1e7d] = 8'hfe; ram[16'h1e7e] = 8'h68; ram[16'h1e7f] = 8'h48; 

ram[16'h1e80] = 8'hc9; ram[16'h1e81] = 8'h30; ram[16'h1e82] = 8'hd0; ram[16'h1e83] = 8'hfe; ram[16'h1e84] = 8'h28; ram[16'h1e85] = 8'ha5; ram[16'h1e86] = 8'h0c; ram[16'h1e87] = 8'hc9; 
ram[16'h1e88] = 8'hfe; ram[16'h1e89] = 8'hd0; ram[16'h1e8a] = 8'hfe; ram[16'h1e8b] = 8'ha9; ram[16'h1e8c] = 8'h01; ram[16'h1e8d] = 8'h85; ram[16'h1e8e] = 8'h0c; ram[16'h1e8f] = 8'ha9; 
ram[16'h1e90] = 8'hff; ram[16'h1e91] = 8'h48; ram[16'h1e92] = 8'ha9; ram[16'h1e93] = 8'h5a; ram[16'h1e94] = 8'h28; ram[16'h1e95] = 8'h07; ram[16'h1e96] = 8'h0c; ram[16'h1e97] = 8'h08; 
ram[16'h1e98] = 8'hc9; ram[16'h1e99] = 8'h5a; ram[16'h1e9a] = 8'hd0; ram[16'h1e9b] = 8'hfe; ram[16'h1e9c] = 8'h68; ram[16'h1e9d] = 8'h48; ram[16'h1e9e] = 8'hc9; ram[16'h1e9f] = 8'hff; 

ram[16'h1ea0] = 8'hd0; ram[16'h1ea1] = 8'hfe; ram[16'h1ea2] = 8'h28; ram[16'h1ea3] = 8'ha5; ram[16'h1ea4] = 8'h0c; ram[16'h1ea5] = 8'hd0; ram[16'h1ea6] = 8'hfe; ram[16'h1ea7] = 8'ha9; 
ram[16'h1ea8] = 8'hff; ram[16'h1ea9] = 8'h85; ram[16'h1eaa] = 8'h0c; ram[16'h1eab] = 8'ha9; ram[16'h1eac] = 8'h00; ram[16'h1ead] = 8'h48; ram[16'h1eae] = 8'ha9; ram[16'h1eaf] = 8'ha5; 
ram[16'h1eb0] = 8'h28; ram[16'h1eb1] = 8'h17; ram[16'h1eb2] = 8'h0c; ram[16'h1eb3] = 8'h08; ram[16'h1eb4] = 8'hc9; ram[16'h1eb5] = 8'ha5; ram[16'h1eb6] = 8'hd0; ram[16'h1eb7] = 8'hfe; 
ram[16'h1eb8] = 8'h68; ram[16'h1eb9] = 8'h48; ram[16'h1eba] = 8'hc9; ram[16'h1ebb] = 8'h30; ram[16'h1ebc] = 8'hd0; ram[16'h1ebd] = 8'hfe; ram[16'h1ebe] = 8'h28; ram[16'h1ebf] = 8'ha5; 

ram[16'h1ec0] = 8'h0c; ram[16'h1ec1] = 8'hc9; ram[16'h1ec2] = 8'hfd; ram[16'h1ec3] = 8'hd0; ram[16'h1ec4] = 8'hfe; ram[16'h1ec5] = 8'ha9; ram[16'h1ec6] = 8'h02; ram[16'h1ec7] = 8'h85; 
ram[16'h1ec8] = 8'h0c; ram[16'h1ec9] = 8'ha9; ram[16'h1eca] = 8'hff; ram[16'h1ecb] = 8'h48; ram[16'h1ecc] = 8'ha9; ram[16'h1ecd] = 8'h5a; ram[16'h1ece] = 8'h28; ram[16'h1ecf] = 8'h17; 
ram[16'h1ed0] = 8'h0c; ram[16'h1ed1] = 8'h08; ram[16'h1ed2] = 8'hc9; ram[16'h1ed3] = 8'h5a; ram[16'h1ed4] = 8'hd0; ram[16'h1ed5] = 8'hfe; ram[16'h1ed6] = 8'h68; ram[16'h1ed7] = 8'h48; 
ram[16'h1ed8] = 8'hc9; ram[16'h1ed9] = 8'hff; ram[16'h1eda] = 8'hd0; ram[16'h1edb] = 8'hfe; ram[16'h1edc] = 8'h28; ram[16'h1edd] = 8'ha5; ram[16'h1ede] = 8'h0c; ram[16'h1edf] = 8'hd0; 

ram[16'h1ee0] = 8'hfe; ram[16'h1ee1] = 8'ha9; ram[16'h1ee2] = 8'hff; ram[16'h1ee3] = 8'h85; ram[16'h1ee4] = 8'h0c; ram[16'h1ee5] = 8'ha9; ram[16'h1ee6] = 8'h00; ram[16'h1ee7] = 8'h48; 
ram[16'h1ee8] = 8'ha9; ram[16'h1ee9] = 8'ha5; ram[16'h1eea] = 8'h28; ram[16'h1eeb] = 8'h27; ram[16'h1eec] = 8'h0c; ram[16'h1eed] = 8'h08; ram[16'h1eee] = 8'hc9; ram[16'h1eef] = 8'ha5; 
ram[16'h1ef0] = 8'hd0; ram[16'h1ef1] = 8'hfe; ram[16'h1ef2] = 8'h68; ram[16'h1ef3] = 8'h48; ram[16'h1ef4] = 8'hc9; ram[16'h1ef5] = 8'h30; ram[16'h1ef6] = 8'hd0; ram[16'h1ef7] = 8'hfe; 
ram[16'h1ef8] = 8'h28; ram[16'h1ef9] = 8'ha5; ram[16'h1efa] = 8'h0c; ram[16'h1efb] = 8'hc9; ram[16'h1efc] = 8'hfb; ram[16'h1efd] = 8'hd0; ram[16'h1efe] = 8'hfe; ram[16'h1eff] = 8'ha9; 

ram[16'h1f00] = 8'h04; ram[16'h1f01] = 8'h85; ram[16'h1f02] = 8'h0c; ram[16'h1f03] = 8'ha9; ram[16'h1f04] = 8'hff; ram[16'h1f05] = 8'h48; ram[16'h1f06] = 8'ha9; ram[16'h1f07] = 8'h5a; 
ram[16'h1f08] = 8'h28; ram[16'h1f09] = 8'h27; ram[16'h1f0a] = 8'h0c; ram[16'h1f0b] = 8'h08; ram[16'h1f0c] = 8'hc9; ram[16'h1f0d] = 8'h5a; ram[16'h1f0e] = 8'hd0; ram[16'h1f0f] = 8'hfe; 
ram[16'h1f10] = 8'h68; ram[16'h1f11] = 8'h48; ram[16'h1f12] = 8'hc9; ram[16'h1f13] = 8'hff; ram[16'h1f14] = 8'hd0; ram[16'h1f15] = 8'hfe; ram[16'h1f16] = 8'h28; ram[16'h1f17] = 8'ha5; 
ram[16'h1f18] = 8'h0c; ram[16'h1f19] = 8'hd0; ram[16'h1f1a] = 8'hfe; ram[16'h1f1b] = 8'ha9; ram[16'h1f1c] = 8'hff; ram[16'h1f1d] = 8'h85; ram[16'h1f1e] = 8'h0c; ram[16'h1f1f] = 8'ha9; 

ram[16'h1f20] = 8'h00; ram[16'h1f21] = 8'h48; ram[16'h1f22] = 8'ha9; ram[16'h1f23] = 8'ha5; ram[16'h1f24] = 8'h28; ram[16'h1f25] = 8'h37; ram[16'h1f26] = 8'h0c; ram[16'h1f27] = 8'h08; 
ram[16'h1f28] = 8'hc9; ram[16'h1f29] = 8'ha5; ram[16'h1f2a] = 8'hd0; ram[16'h1f2b] = 8'hfe; ram[16'h1f2c] = 8'h68; ram[16'h1f2d] = 8'h48; ram[16'h1f2e] = 8'hc9; ram[16'h1f2f] = 8'h30; 
ram[16'h1f30] = 8'hd0; ram[16'h1f31] = 8'hfe; ram[16'h1f32] = 8'h28; ram[16'h1f33] = 8'ha5; ram[16'h1f34] = 8'h0c; ram[16'h1f35] = 8'hc9; ram[16'h1f36] = 8'hf7; ram[16'h1f37] = 8'hd0; 
ram[16'h1f38] = 8'hfe; ram[16'h1f39] = 8'ha9; ram[16'h1f3a] = 8'h08; ram[16'h1f3b] = 8'h85; ram[16'h1f3c] = 8'h0c; ram[16'h1f3d] = 8'ha9; ram[16'h1f3e] = 8'hff; ram[16'h1f3f] = 8'h48; 

ram[16'h1f40] = 8'ha9; ram[16'h1f41] = 8'h5a; ram[16'h1f42] = 8'h28; ram[16'h1f43] = 8'h37; ram[16'h1f44] = 8'h0c; ram[16'h1f45] = 8'h08; ram[16'h1f46] = 8'hc9; ram[16'h1f47] = 8'h5a; 
ram[16'h1f48] = 8'hd0; ram[16'h1f49] = 8'hfe; ram[16'h1f4a] = 8'h68; ram[16'h1f4b] = 8'h48; ram[16'h1f4c] = 8'hc9; ram[16'h1f4d] = 8'hff; ram[16'h1f4e] = 8'hd0; ram[16'h1f4f] = 8'hfe; 
ram[16'h1f50] = 8'h28; ram[16'h1f51] = 8'ha5; ram[16'h1f52] = 8'h0c; ram[16'h1f53] = 8'hd0; ram[16'h1f54] = 8'hfe; ram[16'h1f55] = 8'ha9; ram[16'h1f56] = 8'hff; ram[16'h1f57] = 8'h85; 
ram[16'h1f58] = 8'h0c; ram[16'h1f59] = 8'ha9; ram[16'h1f5a] = 8'h00; ram[16'h1f5b] = 8'h48; ram[16'h1f5c] = 8'ha9; ram[16'h1f5d] = 8'ha5; ram[16'h1f5e] = 8'h28; ram[16'h1f5f] = 8'h47; 

ram[16'h1f60] = 8'h0c; ram[16'h1f61] = 8'h08; ram[16'h1f62] = 8'hc9; ram[16'h1f63] = 8'ha5; ram[16'h1f64] = 8'hd0; ram[16'h1f65] = 8'hfe; ram[16'h1f66] = 8'h68; ram[16'h1f67] = 8'h48; 
ram[16'h1f68] = 8'hc9; ram[16'h1f69] = 8'h30; ram[16'h1f6a] = 8'hd0; ram[16'h1f6b] = 8'hfe; ram[16'h1f6c] = 8'h28; ram[16'h1f6d] = 8'ha5; ram[16'h1f6e] = 8'h0c; ram[16'h1f6f] = 8'hc9; 
ram[16'h1f70] = 8'hef; ram[16'h1f71] = 8'hd0; ram[16'h1f72] = 8'hfe; ram[16'h1f73] = 8'ha9; ram[16'h1f74] = 8'h10; ram[16'h1f75] = 8'h85; ram[16'h1f76] = 8'h0c; ram[16'h1f77] = 8'ha9; 
ram[16'h1f78] = 8'hff; ram[16'h1f79] = 8'h48; ram[16'h1f7a] = 8'ha9; ram[16'h1f7b] = 8'h5a; ram[16'h1f7c] = 8'h28; ram[16'h1f7d] = 8'h47; ram[16'h1f7e] = 8'h0c; ram[16'h1f7f] = 8'h08; 

ram[16'h1f80] = 8'hc9; ram[16'h1f81] = 8'h5a; ram[16'h1f82] = 8'hd0; ram[16'h1f83] = 8'hfe; ram[16'h1f84] = 8'h68; ram[16'h1f85] = 8'h48; ram[16'h1f86] = 8'hc9; ram[16'h1f87] = 8'hff; 
ram[16'h1f88] = 8'hd0; ram[16'h1f89] = 8'hfe; ram[16'h1f8a] = 8'h28; ram[16'h1f8b] = 8'ha5; ram[16'h1f8c] = 8'h0c; ram[16'h1f8d] = 8'hd0; ram[16'h1f8e] = 8'hfe; ram[16'h1f8f] = 8'ha9; 
ram[16'h1f90] = 8'hff; ram[16'h1f91] = 8'h85; ram[16'h1f92] = 8'h0c; ram[16'h1f93] = 8'ha9; ram[16'h1f94] = 8'h00; ram[16'h1f95] = 8'h48; ram[16'h1f96] = 8'ha9; ram[16'h1f97] = 8'ha5; 
ram[16'h1f98] = 8'h28; ram[16'h1f99] = 8'h57; ram[16'h1f9a] = 8'h0c; ram[16'h1f9b] = 8'h08; ram[16'h1f9c] = 8'hc9; ram[16'h1f9d] = 8'ha5; ram[16'h1f9e] = 8'hd0; ram[16'h1f9f] = 8'hfe; 

ram[16'h1fa0] = 8'h68; ram[16'h1fa1] = 8'h48; ram[16'h1fa2] = 8'hc9; ram[16'h1fa3] = 8'h30; ram[16'h1fa4] = 8'hd0; ram[16'h1fa5] = 8'hfe; ram[16'h1fa6] = 8'h28; ram[16'h1fa7] = 8'ha5; 
ram[16'h1fa8] = 8'h0c; ram[16'h1fa9] = 8'hc9; ram[16'h1faa] = 8'hdf; ram[16'h1fab] = 8'hd0; ram[16'h1fac] = 8'hfe; ram[16'h1fad] = 8'ha9; ram[16'h1fae] = 8'h20; ram[16'h1faf] = 8'h85; 
ram[16'h1fb0] = 8'h0c; ram[16'h1fb1] = 8'ha9; ram[16'h1fb2] = 8'hff; ram[16'h1fb3] = 8'h48; ram[16'h1fb4] = 8'ha9; ram[16'h1fb5] = 8'h5a; ram[16'h1fb6] = 8'h28; ram[16'h1fb7] = 8'h57; 
ram[16'h1fb8] = 8'h0c; ram[16'h1fb9] = 8'h08; ram[16'h1fba] = 8'hc9; ram[16'h1fbb] = 8'h5a; ram[16'h1fbc] = 8'hd0; ram[16'h1fbd] = 8'hfe; ram[16'h1fbe] = 8'h68; ram[16'h1fbf] = 8'h48; 

ram[16'h1fc0] = 8'hc9; ram[16'h1fc1] = 8'hff; ram[16'h1fc2] = 8'hd0; ram[16'h1fc3] = 8'hfe; ram[16'h1fc4] = 8'h28; ram[16'h1fc5] = 8'ha5; ram[16'h1fc6] = 8'h0c; ram[16'h1fc7] = 8'hd0; 
ram[16'h1fc8] = 8'hfe; ram[16'h1fc9] = 8'ha9; ram[16'h1fca] = 8'hff; ram[16'h1fcb] = 8'h85; ram[16'h1fcc] = 8'h0c; ram[16'h1fcd] = 8'ha9; ram[16'h1fce] = 8'h00; ram[16'h1fcf] = 8'h48; 
ram[16'h1fd0] = 8'ha9; ram[16'h1fd1] = 8'ha5; ram[16'h1fd2] = 8'h28; ram[16'h1fd3] = 8'h67; ram[16'h1fd4] = 8'h0c; ram[16'h1fd5] = 8'h08; ram[16'h1fd6] = 8'hc9; ram[16'h1fd7] = 8'ha5; 
ram[16'h1fd8] = 8'hd0; ram[16'h1fd9] = 8'hfe; ram[16'h1fda] = 8'h68; ram[16'h1fdb] = 8'h48; ram[16'h1fdc] = 8'hc9; ram[16'h1fdd] = 8'h30; ram[16'h1fde] = 8'hd0; ram[16'h1fdf] = 8'hfe; 

ram[16'h1fe0] = 8'h28; ram[16'h1fe1] = 8'ha5; ram[16'h1fe2] = 8'h0c; ram[16'h1fe3] = 8'hc9; ram[16'h1fe4] = 8'hbf; ram[16'h1fe5] = 8'hd0; ram[16'h1fe6] = 8'hfe; ram[16'h1fe7] = 8'ha9; 
ram[16'h1fe8] = 8'h40; ram[16'h1fe9] = 8'h85; ram[16'h1fea] = 8'h0c; ram[16'h1feb] = 8'ha9; ram[16'h1fec] = 8'hff; ram[16'h1fed] = 8'h48; ram[16'h1fee] = 8'ha9; ram[16'h1fef] = 8'h5a; 
ram[16'h1ff0] = 8'h28; ram[16'h1ff1] = 8'h67; ram[16'h1ff2] = 8'h0c; ram[16'h1ff3] = 8'h08; ram[16'h1ff4] = 8'hc9; ram[16'h1ff5] = 8'h5a; ram[16'h1ff6] = 8'hd0; ram[16'h1ff7] = 8'hfe; 
ram[16'h1ff8] = 8'h68; ram[16'h1ff9] = 8'h48; ram[16'h1ffa] = 8'hc9; ram[16'h1ffb] = 8'hff; ram[16'h1ffc] = 8'hd0; ram[16'h1ffd] = 8'hfe; ram[16'h1ffe] = 8'h28; ram[16'h1fff] = 8'ha5; 

ram[16'h2000] = 8'h0c; ram[16'h2001] = 8'hd0; ram[16'h2002] = 8'hfe; ram[16'h2003] = 8'ha9; ram[16'h2004] = 8'hff; ram[16'h2005] = 8'h85; ram[16'h2006] = 8'h0c; ram[16'h2007] = 8'ha9; 
ram[16'h2008] = 8'h00; ram[16'h2009] = 8'h48; ram[16'h200a] = 8'ha9; ram[16'h200b] = 8'ha5; ram[16'h200c] = 8'h28; ram[16'h200d] = 8'h77; ram[16'h200e] = 8'h0c; ram[16'h200f] = 8'h08; 
ram[16'h2010] = 8'hc9; ram[16'h2011] = 8'ha5; ram[16'h2012] = 8'hd0; ram[16'h2013] = 8'hfe; ram[16'h2014] = 8'h68; ram[16'h2015] = 8'h48; ram[16'h2016] = 8'hc9; ram[16'h2017] = 8'h30; 
ram[16'h2018] = 8'hd0; ram[16'h2019] = 8'hfe; ram[16'h201a] = 8'h28; ram[16'h201b] = 8'ha5; ram[16'h201c] = 8'h0c; ram[16'h201d] = 8'hc9; ram[16'h201e] = 8'h7f; ram[16'h201f] = 8'hd0; 

ram[16'h2020] = 8'hfe; ram[16'h2021] = 8'ha9; ram[16'h2022] = 8'h80; ram[16'h2023] = 8'h85; ram[16'h2024] = 8'h0c; ram[16'h2025] = 8'ha9; ram[16'h2026] = 8'hff; ram[16'h2027] = 8'h48; 
ram[16'h2028] = 8'ha9; ram[16'h2029] = 8'h5a; ram[16'h202a] = 8'h28; ram[16'h202b] = 8'h77; ram[16'h202c] = 8'h0c; ram[16'h202d] = 8'h08; ram[16'h202e] = 8'hc9; ram[16'h202f] = 8'h5a; 
ram[16'h2030] = 8'hd0; ram[16'h2031] = 8'hfe; ram[16'h2032] = 8'h68; ram[16'h2033] = 8'h48; ram[16'h2034] = 8'hc9; ram[16'h2035] = 8'hff; ram[16'h2036] = 8'hd0; ram[16'h2037] = 8'hfe; 
ram[16'h2038] = 8'h28; ram[16'h2039] = 8'ha5; ram[16'h203a] = 8'h0c; ram[16'h203b] = 8'hd0; ram[16'h203c] = 8'hfe; ram[16'h203d] = 8'ha9; ram[16'h203e] = 8'hfe; ram[16'h203f] = 8'h85; 

ram[16'h2040] = 8'h0c; ram[16'h2041] = 8'ha9; ram[16'h2042] = 8'h00; ram[16'h2043] = 8'h48; ram[16'h2044] = 8'ha9; ram[16'h2045] = 8'ha5; ram[16'h2046] = 8'h28; ram[16'h2047] = 8'h87; 
ram[16'h2048] = 8'h0c; ram[16'h2049] = 8'h08; ram[16'h204a] = 8'hc9; ram[16'h204b] = 8'ha5; ram[16'h204c] = 8'hd0; ram[16'h204d] = 8'hfe; ram[16'h204e] = 8'h68; ram[16'h204f] = 8'h48; 
ram[16'h2050] = 8'hc9; ram[16'h2051] = 8'h30; ram[16'h2052] = 8'hd0; ram[16'h2053] = 8'hfe; ram[16'h2054] = 8'h28; ram[16'h2055] = 8'ha5; ram[16'h2056] = 8'h0c; ram[16'h2057] = 8'hc9; 
ram[16'h2058] = 8'hff; ram[16'h2059] = 8'hd0; ram[16'h205a] = 8'hfe; ram[16'h205b] = 8'ha9; ram[16'h205c] = 8'h00; ram[16'h205d] = 8'h85; ram[16'h205e] = 8'h0c; ram[16'h205f] = 8'ha9; 

ram[16'h2060] = 8'hff; ram[16'h2061] = 8'h48; ram[16'h2062] = 8'ha9; ram[16'h2063] = 8'h5a; ram[16'h2064] = 8'h28; ram[16'h2065] = 8'h87; ram[16'h2066] = 8'h0c; ram[16'h2067] = 8'h08; 
ram[16'h2068] = 8'hc9; ram[16'h2069] = 8'h5a; ram[16'h206a] = 8'hd0; ram[16'h206b] = 8'hfe; ram[16'h206c] = 8'h68; ram[16'h206d] = 8'h48; ram[16'h206e] = 8'hc9; ram[16'h206f] = 8'hff; 
ram[16'h2070] = 8'hd0; ram[16'h2071] = 8'hfe; ram[16'h2072] = 8'h28; ram[16'h2073] = 8'ha5; ram[16'h2074] = 8'h0c; ram[16'h2075] = 8'hc9; ram[16'h2076] = 8'h01; ram[16'h2077] = 8'hd0; 
ram[16'h2078] = 8'hfe; ram[16'h2079] = 8'ha9; ram[16'h207a] = 8'hfd; ram[16'h207b] = 8'h85; ram[16'h207c] = 8'h0c; ram[16'h207d] = 8'ha9; ram[16'h207e] = 8'h00; ram[16'h207f] = 8'h48; 

ram[16'h2080] = 8'ha9; ram[16'h2081] = 8'ha5; ram[16'h2082] = 8'h28; ram[16'h2083] = 8'h97; ram[16'h2084] = 8'h0c; ram[16'h2085] = 8'h08; ram[16'h2086] = 8'hc9; ram[16'h2087] = 8'ha5; 
ram[16'h2088] = 8'hd0; ram[16'h2089] = 8'hfe; ram[16'h208a] = 8'h68; ram[16'h208b] = 8'h48; ram[16'h208c] = 8'hc9; ram[16'h208d] = 8'h30; ram[16'h208e] = 8'hd0; ram[16'h208f] = 8'hfe; 
ram[16'h2090] = 8'h28; ram[16'h2091] = 8'ha5; ram[16'h2092] = 8'h0c; ram[16'h2093] = 8'hc9; ram[16'h2094] = 8'hff; ram[16'h2095] = 8'hd0; ram[16'h2096] = 8'hfe; ram[16'h2097] = 8'ha9; 
ram[16'h2098] = 8'h00; ram[16'h2099] = 8'h85; ram[16'h209a] = 8'h0c; ram[16'h209b] = 8'ha9; ram[16'h209c] = 8'hff; ram[16'h209d] = 8'h48; ram[16'h209e] = 8'ha9; ram[16'h209f] = 8'h5a; 

ram[16'h20a0] = 8'h28; ram[16'h20a1] = 8'h97; ram[16'h20a2] = 8'h0c; ram[16'h20a3] = 8'h08; ram[16'h20a4] = 8'hc9; ram[16'h20a5] = 8'h5a; ram[16'h20a6] = 8'hd0; ram[16'h20a7] = 8'hfe; 
ram[16'h20a8] = 8'h68; ram[16'h20a9] = 8'h48; ram[16'h20aa] = 8'hc9; ram[16'h20ab] = 8'hff; ram[16'h20ac] = 8'hd0; ram[16'h20ad] = 8'hfe; ram[16'h20ae] = 8'h28; ram[16'h20af] = 8'ha5; 
ram[16'h20b0] = 8'h0c; ram[16'h20b1] = 8'hc9; ram[16'h20b2] = 8'h02; ram[16'h20b3] = 8'hd0; ram[16'h20b4] = 8'hfe; ram[16'h20b5] = 8'ha9; ram[16'h20b6] = 8'hfb; ram[16'h20b7] = 8'h85; 
ram[16'h20b8] = 8'h0c; ram[16'h20b9] = 8'ha9; ram[16'h20ba] = 8'h00; ram[16'h20bb] = 8'h48; ram[16'h20bc] = 8'ha9; ram[16'h20bd] = 8'ha5; ram[16'h20be] = 8'h28; ram[16'h20bf] = 8'ha7; 

ram[16'h20c0] = 8'h0c; ram[16'h20c1] = 8'h08; ram[16'h20c2] = 8'hc9; ram[16'h20c3] = 8'ha5; ram[16'h20c4] = 8'hd0; ram[16'h20c5] = 8'hfe; ram[16'h20c6] = 8'h68; ram[16'h20c7] = 8'h48; 
ram[16'h20c8] = 8'hc9; ram[16'h20c9] = 8'h30; ram[16'h20ca] = 8'hd0; ram[16'h20cb] = 8'hfe; ram[16'h20cc] = 8'h28; ram[16'h20cd] = 8'ha5; ram[16'h20ce] = 8'h0c; ram[16'h20cf] = 8'hc9; 
ram[16'h20d0] = 8'hff; ram[16'h20d1] = 8'hd0; ram[16'h20d2] = 8'hfe; ram[16'h20d3] = 8'ha9; ram[16'h20d4] = 8'h00; ram[16'h20d5] = 8'h85; ram[16'h20d6] = 8'h0c; ram[16'h20d7] = 8'ha9; 
ram[16'h20d8] = 8'hff; ram[16'h20d9] = 8'h48; ram[16'h20da] = 8'ha9; ram[16'h20db] = 8'h5a; ram[16'h20dc] = 8'h28; ram[16'h20dd] = 8'ha7; ram[16'h20de] = 8'h0c; ram[16'h20df] = 8'h08; 

ram[16'h20e0] = 8'hc9; ram[16'h20e1] = 8'h5a; ram[16'h20e2] = 8'hd0; ram[16'h20e3] = 8'hfe; ram[16'h20e4] = 8'h68; ram[16'h20e5] = 8'h48; ram[16'h20e6] = 8'hc9; ram[16'h20e7] = 8'hff; 
ram[16'h20e8] = 8'hd0; ram[16'h20e9] = 8'hfe; ram[16'h20ea] = 8'h28; ram[16'h20eb] = 8'ha5; ram[16'h20ec] = 8'h0c; ram[16'h20ed] = 8'hc9; ram[16'h20ee] = 8'h04; ram[16'h20ef] = 8'hd0; 
ram[16'h20f0] = 8'hfe; ram[16'h20f1] = 8'ha9; ram[16'h20f2] = 8'hf7; ram[16'h20f3] = 8'h85; ram[16'h20f4] = 8'h0c; ram[16'h20f5] = 8'ha9; ram[16'h20f6] = 8'h00; ram[16'h20f7] = 8'h48; 
ram[16'h20f8] = 8'ha9; ram[16'h20f9] = 8'ha5; ram[16'h20fa] = 8'h28; ram[16'h20fb] = 8'hb7; ram[16'h20fc] = 8'h0c; ram[16'h20fd] = 8'h08; ram[16'h20fe] = 8'hc9; ram[16'h20ff] = 8'ha5; 

ram[16'h2100] = 8'hd0; ram[16'h2101] = 8'hfe; ram[16'h2102] = 8'h68; ram[16'h2103] = 8'h48; ram[16'h2104] = 8'hc9; ram[16'h2105] = 8'h30; ram[16'h2106] = 8'hd0; ram[16'h2107] = 8'hfe; 
ram[16'h2108] = 8'h28; ram[16'h2109] = 8'ha5; ram[16'h210a] = 8'h0c; ram[16'h210b] = 8'hc9; ram[16'h210c] = 8'hff; ram[16'h210d] = 8'hd0; ram[16'h210e] = 8'hfe; ram[16'h210f] = 8'ha9; 
ram[16'h2110] = 8'h00; ram[16'h2111] = 8'h85; ram[16'h2112] = 8'h0c; ram[16'h2113] = 8'ha9; ram[16'h2114] = 8'hff; ram[16'h2115] = 8'h48; ram[16'h2116] = 8'ha9; ram[16'h2117] = 8'h5a; 
ram[16'h2118] = 8'h28; ram[16'h2119] = 8'hb7; ram[16'h211a] = 8'h0c; ram[16'h211b] = 8'h08; ram[16'h211c] = 8'hc9; ram[16'h211d] = 8'h5a; ram[16'h211e] = 8'hd0; ram[16'h211f] = 8'hfe; 

ram[16'h2120] = 8'h68; ram[16'h2121] = 8'h48; ram[16'h2122] = 8'hc9; ram[16'h2123] = 8'hff; ram[16'h2124] = 8'hd0; ram[16'h2125] = 8'hfe; ram[16'h2126] = 8'h28; ram[16'h2127] = 8'ha5; 
ram[16'h2128] = 8'h0c; ram[16'h2129] = 8'hc9; ram[16'h212a] = 8'h08; ram[16'h212b] = 8'hd0; ram[16'h212c] = 8'hfe; ram[16'h212d] = 8'ha9; ram[16'h212e] = 8'hef; ram[16'h212f] = 8'h85; 
ram[16'h2130] = 8'h0c; ram[16'h2131] = 8'ha9; ram[16'h2132] = 8'h00; ram[16'h2133] = 8'h48; ram[16'h2134] = 8'ha9; ram[16'h2135] = 8'ha5; ram[16'h2136] = 8'h28; ram[16'h2137] = 8'hc7; 
ram[16'h2138] = 8'h0c; ram[16'h2139] = 8'h08; ram[16'h213a] = 8'hc9; ram[16'h213b] = 8'ha5; ram[16'h213c] = 8'hd0; ram[16'h213d] = 8'hfe; ram[16'h213e] = 8'h68; ram[16'h213f] = 8'h48; 

ram[16'h2140] = 8'hc9; ram[16'h2141] = 8'h30; ram[16'h2142] = 8'hd0; ram[16'h2143] = 8'hfe; ram[16'h2144] = 8'h28; ram[16'h2145] = 8'ha5; ram[16'h2146] = 8'h0c; ram[16'h2147] = 8'hc9; 
ram[16'h2148] = 8'hff; ram[16'h2149] = 8'hd0; ram[16'h214a] = 8'hfe; ram[16'h214b] = 8'ha9; ram[16'h214c] = 8'h00; ram[16'h214d] = 8'h85; ram[16'h214e] = 8'h0c; ram[16'h214f] = 8'ha9; 
ram[16'h2150] = 8'hff; ram[16'h2151] = 8'h48; ram[16'h2152] = 8'ha9; ram[16'h2153] = 8'h5a; ram[16'h2154] = 8'h28; ram[16'h2155] = 8'hc7; ram[16'h2156] = 8'h0c; ram[16'h2157] = 8'h08; 
ram[16'h2158] = 8'hc9; ram[16'h2159] = 8'h5a; ram[16'h215a] = 8'hd0; ram[16'h215b] = 8'hfe; ram[16'h215c] = 8'h68; ram[16'h215d] = 8'h48; ram[16'h215e] = 8'hc9; ram[16'h215f] = 8'hff; 

ram[16'h2160] = 8'hd0; ram[16'h2161] = 8'hfe; ram[16'h2162] = 8'h28; ram[16'h2163] = 8'ha5; ram[16'h2164] = 8'h0c; ram[16'h2165] = 8'hc9; ram[16'h2166] = 8'h10; ram[16'h2167] = 8'hd0; 
ram[16'h2168] = 8'hfe; ram[16'h2169] = 8'ha9; ram[16'h216a] = 8'hdf; ram[16'h216b] = 8'h85; ram[16'h216c] = 8'h0c; ram[16'h216d] = 8'ha9; ram[16'h216e] = 8'h00; ram[16'h216f] = 8'h48; 
ram[16'h2170] = 8'ha9; ram[16'h2171] = 8'ha5; ram[16'h2172] = 8'h28; ram[16'h2173] = 8'hd7; ram[16'h2174] = 8'h0c; ram[16'h2175] = 8'h08; ram[16'h2176] = 8'hc9; ram[16'h2177] = 8'ha5; 
ram[16'h2178] = 8'hd0; ram[16'h2179] = 8'hfe; ram[16'h217a] = 8'h68; ram[16'h217b] = 8'h48; ram[16'h217c] = 8'hc9; ram[16'h217d] = 8'h30; ram[16'h217e] = 8'hd0; ram[16'h217f] = 8'hfe; 

ram[16'h2180] = 8'h28; ram[16'h2181] = 8'ha5; ram[16'h2182] = 8'h0c; ram[16'h2183] = 8'hc9; ram[16'h2184] = 8'hff; ram[16'h2185] = 8'hd0; ram[16'h2186] = 8'hfe; ram[16'h2187] = 8'ha9; 
ram[16'h2188] = 8'h00; ram[16'h2189] = 8'h85; ram[16'h218a] = 8'h0c; ram[16'h218b] = 8'ha9; ram[16'h218c] = 8'hff; ram[16'h218d] = 8'h48; ram[16'h218e] = 8'ha9; ram[16'h218f] = 8'h5a; 
ram[16'h2190] = 8'h28; ram[16'h2191] = 8'hd7; ram[16'h2192] = 8'h0c; ram[16'h2193] = 8'h08; ram[16'h2194] = 8'hc9; ram[16'h2195] = 8'h5a; ram[16'h2196] = 8'hd0; ram[16'h2197] = 8'hfe; 
ram[16'h2198] = 8'h68; ram[16'h2199] = 8'h48; ram[16'h219a] = 8'hc9; ram[16'h219b] = 8'hff; ram[16'h219c] = 8'hd0; ram[16'h219d] = 8'hfe; ram[16'h219e] = 8'h28; ram[16'h219f] = 8'ha5; 

ram[16'h21a0] = 8'h0c; ram[16'h21a1] = 8'hc9; ram[16'h21a2] = 8'h20; ram[16'h21a3] = 8'hd0; ram[16'h21a4] = 8'hfe; ram[16'h21a5] = 8'ha9; ram[16'h21a6] = 8'hbf; ram[16'h21a7] = 8'h85; 
ram[16'h21a8] = 8'h0c; ram[16'h21a9] = 8'ha9; ram[16'h21aa] = 8'h00; ram[16'h21ab] = 8'h48; ram[16'h21ac] = 8'ha9; ram[16'h21ad] = 8'ha5; ram[16'h21ae] = 8'h28; ram[16'h21af] = 8'he7; 
ram[16'h21b0] = 8'h0c; ram[16'h21b1] = 8'h08; ram[16'h21b2] = 8'hc9; ram[16'h21b3] = 8'ha5; ram[16'h21b4] = 8'hd0; ram[16'h21b5] = 8'hfe; ram[16'h21b6] = 8'h68; ram[16'h21b7] = 8'h48; 
ram[16'h21b8] = 8'hc9; ram[16'h21b9] = 8'h30; ram[16'h21ba] = 8'hd0; ram[16'h21bb] = 8'hfe; ram[16'h21bc] = 8'h28; ram[16'h21bd] = 8'ha5; ram[16'h21be] = 8'h0c; ram[16'h21bf] = 8'hc9; 

ram[16'h21c0] = 8'hff; ram[16'h21c1] = 8'hd0; ram[16'h21c2] = 8'hfe; ram[16'h21c3] = 8'ha9; ram[16'h21c4] = 8'h00; ram[16'h21c5] = 8'h85; ram[16'h21c6] = 8'h0c; ram[16'h21c7] = 8'ha9; 
ram[16'h21c8] = 8'hff; ram[16'h21c9] = 8'h48; ram[16'h21ca] = 8'ha9; ram[16'h21cb] = 8'h5a; ram[16'h21cc] = 8'h28; ram[16'h21cd] = 8'he7; ram[16'h21ce] = 8'h0c; ram[16'h21cf] = 8'h08; 
ram[16'h21d0] = 8'hc9; ram[16'h21d1] = 8'h5a; ram[16'h21d2] = 8'hd0; ram[16'h21d3] = 8'hfe; ram[16'h21d4] = 8'h68; ram[16'h21d5] = 8'h48; ram[16'h21d6] = 8'hc9; ram[16'h21d7] = 8'hff; 
ram[16'h21d8] = 8'hd0; ram[16'h21d9] = 8'hfe; ram[16'h21da] = 8'h28; ram[16'h21db] = 8'ha5; ram[16'h21dc] = 8'h0c; ram[16'h21dd] = 8'hc9; ram[16'h21de] = 8'h40; ram[16'h21df] = 8'hd0; 

ram[16'h21e0] = 8'hfe; ram[16'h21e1] = 8'ha9; ram[16'h21e2] = 8'h7f; ram[16'h21e3] = 8'h85; ram[16'h21e4] = 8'h0c; ram[16'h21e5] = 8'ha9; ram[16'h21e6] = 8'h00; ram[16'h21e7] = 8'h48; 
ram[16'h21e8] = 8'ha9; ram[16'h21e9] = 8'ha5; ram[16'h21ea] = 8'h28; ram[16'h21eb] = 8'hf7; ram[16'h21ec] = 8'h0c; ram[16'h21ed] = 8'h08; ram[16'h21ee] = 8'hc9; ram[16'h21ef] = 8'ha5; 
ram[16'h21f0] = 8'hd0; ram[16'h21f1] = 8'hfe; ram[16'h21f2] = 8'h68; ram[16'h21f3] = 8'h48; ram[16'h21f4] = 8'hc9; ram[16'h21f5] = 8'h30; ram[16'h21f6] = 8'hd0; ram[16'h21f7] = 8'hfe; 
ram[16'h21f8] = 8'h28; ram[16'h21f9] = 8'ha5; ram[16'h21fa] = 8'h0c; ram[16'h21fb] = 8'hc9; ram[16'h21fc] = 8'hff; ram[16'h21fd] = 8'hd0; ram[16'h21fe] = 8'hfe; ram[16'h21ff] = 8'ha9; 

ram[16'h2200] = 8'h00; ram[16'h2201] = 8'h85; ram[16'h2202] = 8'h0c; ram[16'h2203] = 8'ha9; ram[16'h2204] = 8'hff; ram[16'h2205] = 8'h48; ram[16'h2206] = 8'ha9; ram[16'h2207] = 8'h5a; 
ram[16'h2208] = 8'h28; ram[16'h2209] = 8'hf7; ram[16'h220a] = 8'h0c; ram[16'h220b] = 8'h08; ram[16'h220c] = 8'hc9; ram[16'h220d] = 8'h5a; ram[16'h220e] = 8'hd0; ram[16'h220f] = 8'hfe; 
ram[16'h2210] = 8'h68; ram[16'h2211] = 8'h48; ram[16'h2212] = 8'hc9; ram[16'h2213] = 8'hff; ram[16'h2214] = 8'hd0; ram[16'h2215] = 8'hfe; ram[16'h2216] = 8'h28; ram[16'h2217] = 8'ha5; 
ram[16'h2218] = 8'h0c; ram[16'h2219] = 8'hc9; ram[16'h221a] = 8'h80; ram[16'h221b] = 8'hd0; ram[16'h221c] = 8'hfe; ram[16'h221d] = 8'he0; ram[16'h221e] = 8'hba; ram[16'h221f] = 8'hd0; 

ram[16'h2220] = 8'hfe; ram[16'h2221] = 8'hc0; ram[16'h2222] = 8'hd0; ram[16'h2223] = 8'hd0; ram[16'h2224] = 8'hfe; ram[16'h2225] = 8'hba; ram[16'h2226] = 8'he0; ram[16'h2227] = 8'hff; 
ram[16'h2228] = 8'hd0; ram[16'h2229] = 8'hfe; ram[16'h222a] = 8'had; ram[16'h222b] = 8'h02; ram[16'h222c] = 8'h02; ram[16'h222d] = 8'hc9; ram[16'h222e] = 8'h11; ram[16'h222f] = 8'hd0; 
ram[16'h2230] = 8'hfe; ram[16'h2231] = 8'ha9; ram[16'h2232] = 8'h12; ram[16'h2233] = 8'h8d; ram[16'h2234] = 8'h02; ram[16'h2235] = 8'h02; ram[16'h2236] = 8'ha2; ram[16'h2237] = 8'hde; 
ram[16'h2238] = 8'ha0; ram[16'h2239] = 8'had; ram[16'h223a] = 8'ha9; ram[16'h223b] = 8'h00; ram[16'h223c] = 8'h48; ram[16'h223d] = 8'ha9; ram[16'h223e] = 8'h80; ram[16'h223f] = 8'h28; 

ram[16'h2240] = 8'hd2; ram[16'h2241] = 8'h2c; ram[16'h2242] = 8'h08; ram[16'h2243] = 8'hc9; ram[16'h2244] = 8'h80; ram[16'h2245] = 8'hd0; ram[16'h2246] = 8'hfe; ram[16'h2247] = 8'h68; 
ram[16'h2248] = 8'h48; ram[16'h2249] = 8'hc9; ram[16'h224a] = 8'h31; ram[16'h224b] = 8'hd0; ram[16'h224c] = 8'hfe; ram[16'h224d] = 8'h28; ram[16'h224e] = 8'ha9; ram[16'h224f] = 8'h00; 
ram[16'h2250] = 8'h48; ram[16'h2251] = 8'ha9; ram[16'h2252] = 8'h7f; ram[16'h2253] = 8'h28; ram[16'h2254] = 8'hd2; ram[16'h2255] = 8'h2c; ram[16'h2256] = 8'h08; ram[16'h2257] = 8'hc9; 
ram[16'h2258] = 8'h7f; ram[16'h2259] = 8'hd0; ram[16'h225a] = 8'hfe; ram[16'h225b] = 8'h68; ram[16'h225c] = 8'h48; ram[16'h225d] = 8'hc9; ram[16'h225e] = 8'h33; ram[16'h225f] = 8'hd0; 

ram[16'h2260] = 8'hfe; ram[16'h2261] = 8'h28; ram[16'h2262] = 8'ha9; ram[16'h2263] = 8'h00; ram[16'h2264] = 8'h48; ram[16'h2265] = 8'ha9; ram[16'h2266] = 8'h7e; ram[16'h2267] = 8'h28; 
ram[16'h2268] = 8'hd2; ram[16'h2269] = 8'h2c; ram[16'h226a] = 8'h08; ram[16'h226b] = 8'hc9; ram[16'h226c] = 8'h7e; ram[16'h226d] = 8'hd0; ram[16'h226e] = 8'hfe; ram[16'h226f] = 8'h68; 
ram[16'h2270] = 8'h48; ram[16'h2271] = 8'hc9; ram[16'h2272] = 8'hb0; ram[16'h2273] = 8'hd0; ram[16'h2274] = 8'hfe; ram[16'h2275] = 8'h28; ram[16'h2276] = 8'ha9; ram[16'h2277] = 8'hff; 
ram[16'h2278] = 8'h48; ram[16'h2279] = 8'ha9; ram[16'h227a] = 8'h80; ram[16'h227b] = 8'h28; ram[16'h227c] = 8'hd2; ram[16'h227d] = 8'h2c; ram[16'h227e] = 8'h08; ram[16'h227f] = 8'hc9; 

ram[16'h2280] = 8'h80; ram[16'h2281] = 8'hd0; ram[16'h2282] = 8'hfe; ram[16'h2283] = 8'h68; ram[16'h2284] = 8'h48; ram[16'h2285] = 8'hc9; ram[16'h2286] = 8'h7d; ram[16'h2287] = 8'hd0; 
ram[16'h2288] = 8'hfe; ram[16'h2289] = 8'h28; ram[16'h228a] = 8'ha9; ram[16'h228b] = 8'hff; ram[16'h228c] = 8'h48; ram[16'h228d] = 8'ha9; ram[16'h228e] = 8'h7f; ram[16'h228f] = 8'h28; 
ram[16'h2290] = 8'hd2; ram[16'h2291] = 8'h2c; ram[16'h2292] = 8'h08; ram[16'h2293] = 8'hc9; ram[16'h2294] = 8'h7f; ram[16'h2295] = 8'hd0; ram[16'h2296] = 8'hfe; ram[16'h2297] = 8'h68; 
ram[16'h2298] = 8'h48; ram[16'h2299] = 8'hc9; ram[16'h229a] = 8'h7f; ram[16'h229b] = 8'hd0; ram[16'h229c] = 8'hfe; ram[16'h229d] = 8'h28; ram[16'h229e] = 8'ha9; ram[16'h229f] = 8'hff; 

ram[16'h22a0] = 8'h48; ram[16'h22a1] = 8'ha9; ram[16'h22a2] = 8'h7e; ram[16'h22a3] = 8'h28; ram[16'h22a4] = 8'hd2; ram[16'h22a5] = 8'h2c; ram[16'h22a6] = 8'h08; ram[16'h22a7] = 8'hc9; 
ram[16'h22a8] = 8'h7e; ram[16'h22a9] = 8'hd0; ram[16'h22aa] = 8'hfe; ram[16'h22ab] = 8'h68; ram[16'h22ac] = 8'h48; ram[16'h22ad] = 8'hc9; ram[16'h22ae] = 8'hfc; ram[16'h22af] = 8'hd0; 
ram[16'h22b0] = 8'hfe; ram[16'h22b1] = 8'h28; ram[16'h22b2] = 8'he0; ram[16'h22b3] = 8'hde; ram[16'h22b4] = 8'hd0; ram[16'h22b5] = 8'hfe; ram[16'h22b6] = 8'hc0; ram[16'h22b7] = 8'had; 
ram[16'h22b8] = 8'hd0; ram[16'h22b9] = 8'hfe; ram[16'h22ba] = 8'hba; ram[16'h22bb] = 8'he0; ram[16'h22bc] = 8'hff; ram[16'h22bd] = 8'hd0; ram[16'h22be] = 8'hfe; ram[16'h22bf] = 8'had; 

ram[16'h22c0] = 8'h02; ram[16'h22c1] = 8'h02; ram[16'h22c2] = 8'hc9; ram[16'h22c3] = 8'h12; ram[16'h22c4] = 8'hd0; ram[16'h22c5] = 8'hfe; ram[16'h22c6] = 8'ha9; ram[16'h22c7] = 8'h13; 
ram[16'h22c8] = 8'h8d; ram[16'h22c9] = 8'h02; ram[16'h22ca] = 8'h02; ram[16'h22cb] = 8'ha2; ram[16'h22cc] = 8'h42; ram[16'h22cd] = 8'ha0; ram[16'h22ce] = 8'h00; ram[16'h22cf] = 8'ha5; 
ram[16'h22d0] = 8'h3a; ram[16'h22d1] = 8'h85; ram[16'h22d2] = 8'h0c; ram[16'h22d3] = 8'ha5; ram[16'h22d4] = 8'h3b; ram[16'h22d5] = 8'h85; ram[16'h22d6] = 8'h0d; ram[16'h22d7] = 8'ha9; 
ram[16'h22d8] = 8'h00; ram[16'h22d9] = 8'h48; ram[16'h22da] = 8'hb9; ram[16'h22db] = 8'h53; ram[16'h22dc] = 8'h02; ram[16'h22dd] = 8'h28; ram[16'h22de] = 8'h32; ram[16'h22df] = 8'h0c; 

ram[16'h22e0] = 8'h08; ram[16'h22e1] = 8'hd9; ram[16'h22e2] = 8'h5b; ram[16'h22e3] = 8'h02; ram[16'h22e4] = 8'hd0; ram[16'h22e5] = 8'hfe; ram[16'h22e6] = 8'h68; ram[16'h22e7] = 8'h49; 
ram[16'h22e8] = 8'h30; ram[16'h22e9] = 8'hd9; ram[16'h22ea] = 8'h5f; ram[16'h22eb] = 8'h02; ram[16'h22ec] = 8'hd0; ram[16'h22ed] = 8'hfe; ram[16'h22ee] = 8'he6; ram[16'h22ef] = 8'h0c; 
ram[16'h22f0] = 8'hc8; ram[16'h22f1] = 8'hc0; ram[16'h22f2] = 8'h04; ram[16'h22f3] = 8'hd0; ram[16'h22f4] = 8'he2; ram[16'h22f5] = 8'h88; ram[16'h22f6] = 8'hc6; ram[16'h22f7] = 8'h0c; 
ram[16'h22f8] = 8'ha9; ram[16'h22f9] = 8'hff; ram[16'h22fa] = 8'h48; ram[16'h22fb] = 8'hb9; ram[16'h22fc] = 8'h53; ram[16'h22fd] = 8'h02; ram[16'h22fe] = 8'h28; ram[16'h22ff] = 8'h32; 

ram[16'h2300] = 8'h0c; ram[16'h2301] = 8'h08; ram[16'h2302] = 8'hd9; ram[16'h2303] = 8'h5b; ram[16'h2304] = 8'h02; ram[16'h2305] = 8'hd0; ram[16'h2306] = 8'hfe; ram[16'h2307] = 8'h68; 
ram[16'h2308] = 8'h49; ram[16'h2309] = 8'h7d; ram[16'h230a] = 8'hd9; ram[16'h230b] = 8'h5f; ram[16'h230c] = 8'h02; ram[16'h230d] = 8'hd0; ram[16'h230e] = 8'hfe; ram[16'h230f] = 8'hc6; 
ram[16'h2310] = 8'h0c; ram[16'h2311] = 8'h88; ram[16'h2312] = 8'h10; ram[16'h2313] = 8'he4; ram[16'h2314] = 8'ha0; ram[16'h2315] = 8'h00; ram[16'h2316] = 8'ha5; ram[16'h2317] = 8'h42; 
ram[16'h2318] = 8'h85; ram[16'h2319] = 8'h0c; ram[16'h231a] = 8'ha5; ram[16'h231b] = 8'h43; ram[16'h231c] = 8'h85; ram[16'h231d] = 8'h0d; ram[16'h231e] = 8'ha9; ram[16'h231f] = 8'h00; 

ram[16'h2320] = 8'h48; ram[16'h2321] = 8'hb9; ram[16'h2322] = 8'h57; ram[16'h2323] = 8'h02; ram[16'h2324] = 8'h28; ram[16'h2325] = 8'h52; ram[16'h2326] = 8'h0c; ram[16'h2327] = 8'h08; 
ram[16'h2328] = 8'hd9; ram[16'h2329] = 8'h5b; ram[16'h232a] = 8'h02; ram[16'h232b] = 8'hd0; ram[16'h232c] = 8'hfe; ram[16'h232d] = 8'h68; ram[16'h232e] = 8'h49; ram[16'h232f] = 8'h30; 
ram[16'h2330] = 8'hd9; ram[16'h2331] = 8'h5f; ram[16'h2332] = 8'h02; ram[16'h2333] = 8'hd0; ram[16'h2334] = 8'hfe; ram[16'h2335] = 8'he6; ram[16'h2336] = 8'h0c; ram[16'h2337] = 8'hc8; 
ram[16'h2338] = 8'hc0; ram[16'h2339] = 8'h04; ram[16'h233a] = 8'hd0; ram[16'h233b] = 8'he2; ram[16'h233c] = 8'h88; ram[16'h233d] = 8'hc6; ram[16'h233e] = 8'h0c; ram[16'h233f] = 8'ha9; 

ram[16'h2340] = 8'hff; ram[16'h2341] = 8'h48; ram[16'h2342] = 8'hb9; ram[16'h2343] = 8'h57; ram[16'h2344] = 8'h02; ram[16'h2345] = 8'h28; ram[16'h2346] = 8'h52; ram[16'h2347] = 8'h0c; 
ram[16'h2348] = 8'h08; ram[16'h2349] = 8'hd9; ram[16'h234a] = 8'h5b; ram[16'h234b] = 8'h02; ram[16'h234c] = 8'hd0; ram[16'h234d] = 8'hfe; ram[16'h234e] = 8'h68; ram[16'h234f] = 8'h49; 
ram[16'h2350] = 8'h7d; ram[16'h2351] = 8'hd9; ram[16'h2352] = 8'h5f; ram[16'h2353] = 8'h02; ram[16'h2354] = 8'hd0; ram[16'h2355] = 8'hfe; ram[16'h2356] = 8'hc6; ram[16'h2357] = 8'h0c; 
ram[16'h2358] = 8'h88; ram[16'h2359] = 8'h10; ram[16'h235a] = 8'he4; ram[16'h235b] = 8'ha0; ram[16'h235c] = 8'h00; ram[16'h235d] = 8'ha5; ram[16'h235e] = 8'h4a; ram[16'h235f] = 8'h85; 

ram[16'h2360] = 8'h0c; ram[16'h2361] = 8'ha5; ram[16'h2362] = 8'h4b; ram[16'h2363] = 8'h85; ram[16'h2364] = 8'h0d; ram[16'h2365] = 8'ha9; ram[16'h2366] = 8'h00; ram[16'h2367] = 8'h48; 
ram[16'h2368] = 8'hb9; ram[16'h2369] = 8'h4f; ram[16'h236a] = 8'h02; ram[16'h236b] = 8'h28; ram[16'h236c] = 8'h12; ram[16'h236d] = 8'h0c; ram[16'h236e] = 8'h08; ram[16'h236f] = 8'hd9; 
ram[16'h2370] = 8'h5b; ram[16'h2371] = 8'h02; ram[16'h2372] = 8'hd0; ram[16'h2373] = 8'hfe; ram[16'h2374] = 8'h68; ram[16'h2375] = 8'h49; ram[16'h2376] = 8'h30; ram[16'h2377] = 8'hd9; 
ram[16'h2378] = 8'h5f; ram[16'h2379] = 8'h02; ram[16'h237a] = 8'hd0; ram[16'h237b] = 8'hfe; ram[16'h237c] = 8'he6; ram[16'h237d] = 8'h0c; ram[16'h237e] = 8'hc8; ram[16'h237f] = 8'hc0; 

ram[16'h2380] = 8'h04; ram[16'h2381] = 8'hd0; ram[16'h2382] = 8'he2; ram[16'h2383] = 8'h88; ram[16'h2384] = 8'hc6; ram[16'h2385] = 8'h0c; ram[16'h2386] = 8'ha9; ram[16'h2387] = 8'hff; 
ram[16'h2388] = 8'h48; ram[16'h2389] = 8'hb9; ram[16'h238a] = 8'h4f; ram[16'h238b] = 8'h02; ram[16'h238c] = 8'h28; ram[16'h238d] = 8'h12; ram[16'h238e] = 8'h0c; ram[16'h238f] = 8'h08; 
ram[16'h2390] = 8'hd9; ram[16'h2391] = 8'h5b; ram[16'h2392] = 8'h02; ram[16'h2393] = 8'hd0; ram[16'h2394] = 8'hfe; ram[16'h2395] = 8'h68; ram[16'h2396] = 8'h49; ram[16'h2397] = 8'h7d; 
ram[16'h2398] = 8'hd9; ram[16'h2399] = 8'h5f; ram[16'h239a] = 8'h02; ram[16'h239b] = 8'hd0; ram[16'h239c] = 8'hfe; ram[16'h239d] = 8'hc6; ram[16'h239e] = 8'h0c; ram[16'h239f] = 8'h88; 

ram[16'h23a0] = 8'h10; ram[16'h23a1] = 8'he4; ram[16'h23a2] = 8'he0; ram[16'h23a3] = 8'h42; ram[16'h23a4] = 8'hd0; ram[16'h23a5] = 8'hfe; ram[16'h23a6] = 8'hba; ram[16'h23a7] = 8'he0; 
ram[16'h23a8] = 8'hff; ram[16'h23a9] = 8'hd0; ram[16'h23aa] = 8'hfe; ram[16'h23ab] = 8'had; ram[16'h23ac] = 8'h02; ram[16'h23ad] = 8'h02; ram[16'h23ae] = 8'hc9; ram[16'h23af] = 8'h13; 
ram[16'h23b0] = 8'hd0; ram[16'h23b1] = 8'hfe; ram[16'h23b2] = 8'ha9; ram[16'h23b3] = 8'h14; ram[16'h23b4] = 8'h8d; ram[16'h23b5] = 8'h02; ram[16'h23b6] = 8'h02; ram[16'h23b7] = 8'h58; 
ram[16'h23b8] = 8'hd8; ram[16'h23b9] = 8'ha2; ram[16'h23ba] = 8'h0e; ram[16'h23bb] = 8'ha0; ram[16'h23bc] = 8'hff; ram[16'h23bd] = 8'ha9; ram[16'h23be] = 8'h00; ram[16'h23bf] = 8'h85; 

ram[16'h23c0] = 8'h0c; ram[16'h23c1] = 8'h85; ram[16'h23c2] = 8'h0d; ram[16'h23c3] = 8'h85; ram[16'h23c4] = 8'h0e; ram[16'h23c5] = 8'h8d; ram[16'h23c6] = 8'h05; ram[16'h23c7] = 8'h02; 
ram[16'h23c8] = 8'h85; ram[16'h23c9] = 8'h0f; ram[16'h23ca] = 8'h85; ram[16'h23cb] = 8'h10; ram[16'h23cc] = 8'ha9; ram[16'h23cd] = 8'hff; ram[16'h23ce] = 8'h85; ram[16'h23cf] = 8'h12; 
ram[16'h23d0] = 8'h8d; ram[16'h23d1] = 8'h06; ram[16'h23d2] = 8'h02; ram[16'h23d3] = 8'ha9; ram[16'h23d4] = 8'h02; ram[16'h23d5] = 8'h85; ram[16'h23d6] = 8'h11; ram[16'h23d7] = 8'h18; 
ram[16'h23d8] = 8'h20; ram[16'h23d9] = 8'h4e; ram[16'h23da] = 8'h26; ram[16'h23db] = 8'he6; ram[16'h23dc] = 8'h0c; ram[16'h23dd] = 8'he6; ram[16'h23de] = 8'h0f; ram[16'h23df] = 8'h08; 

ram[16'h23e0] = 8'h08; ram[16'h23e1] = 8'h68; ram[16'h23e2] = 8'h29; ram[16'h23e3] = 8'h82; ram[16'h23e4] = 8'h28; ram[16'h23e5] = 8'hd0; ram[16'h23e6] = 8'h02; ram[16'h23e7] = 8'he6; 
ram[16'h23e8] = 8'h10; ram[16'h23e9] = 8'h05; ram[16'h23ea] = 8'h10; ram[16'h23eb] = 8'h85; ram[16'h23ec] = 8'h11; ram[16'h23ed] = 8'h38; ram[16'h23ee] = 8'h20; ram[16'h23ef] = 8'h4e; 
ram[16'h23f0] = 8'h26; ram[16'h23f1] = 8'hc6; ram[16'h23f2] = 8'h0c; ram[16'h23f3] = 8'he6; ram[16'h23f4] = 8'h0d; ram[16'h23f5] = 8'hd0; ram[16'h23f6] = 8'he0; ram[16'h23f7] = 8'ha9; 
ram[16'h23f8] = 8'h00; ram[16'h23f9] = 8'h85; ram[16'h23fa] = 8'h10; ram[16'h23fb] = 8'hee; ram[16'h23fc] = 8'h05; ram[16'h23fd] = 8'h02; ram[16'h23fe] = 8'he6; ram[16'h23ff] = 8'h0e; 

ram[16'h2400] = 8'h08; ram[16'h2401] = 8'h68; ram[16'h2402] = 8'h29; ram[16'h2403] = 8'h82; ram[16'h2404] = 8'h85; ram[16'h2405] = 8'h11; ram[16'h2406] = 8'hc6; ram[16'h2407] = 8'h12; 
ram[16'h2408] = 8'hce; ram[16'h2409] = 8'h06; ram[16'h240a] = 8'h02; ram[16'h240b] = 8'ha5; ram[16'h240c] = 8'h0e; ram[16'h240d] = 8'h85; ram[16'h240e] = 8'h0f; ram[16'h240f] = 8'hd0; 
ram[16'h2410] = 8'hc6; ram[16'h2411] = 8'he0; ram[16'h2412] = 8'h0e; ram[16'h2413] = 8'hd0; ram[16'h2414] = 8'hfe; ram[16'h2415] = 8'hc0; ram[16'h2416] = 8'hff; ram[16'h2417] = 8'hd0; 
ram[16'h2418] = 8'hfe; ram[16'h2419] = 8'hba; ram[16'h241a] = 8'he0; ram[16'h241b] = 8'hff; ram[16'h241c] = 8'hd0; ram[16'h241d] = 8'hfe; ram[16'h241e] = 8'had; ram[16'h241f] = 8'h02; 

ram[16'h2420] = 8'h02; ram[16'h2421] = 8'hc9; ram[16'h2422] = 8'h14; ram[16'h2423] = 8'hd0; ram[16'h2424] = 8'hfe; ram[16'h2425] = 8'ha9; ram[16'h2426] = 8'h15; ram[16'h2427] = 8'h8d; 
ram[16'h2428] = 8'h02; ram[16'h2429] = 8'h02; ram[16'h242a] = 8'hf8; ram[16'h242b] = 8'ha2; ram[16'h242c] = 8'h0e; ram[16'h242d] = 8'ha0; ram[16'h242e] = 8'hff; ram[16'h242f] = 8'ha9; 
ram[16'h2430] = 8'h99; ram[16'h2431] = 8'h85; ram[16'h2432] = 8'h0d; ram[16'h2433] = 8'h85; ram[16'h2434] = 8'h0e; ram[16'h2435] = 8'h8d; ram[16'h2436] = 8'h05; ram[16'h2437] = 8'h02; 
ram[16'h2438] = 8'h85; ram[16'h2439] = 8'h0f; ram[16'h243a] = 8'ha9; ram[16'h243b] = 8'h01; ram[16'h243c] = 8'h85; ram[16'h243d] = 8'h0c; ram[16'h243e] = 8'h85; ram[16'h243f] = 8'h10; 

ram[16'h2440] = 8'ha9; ram[16'h2441] = 8'h81; ram[16'h2442] = 8'h85; ram[16'h2443] = 8'h11; ram[16'h2444] = 8'ha9; ram[16'h2445] = 8'h00; ram[16'h2446] = 8'h85; ram[16'h2447] = 8'h12; 
ram[16'h2448] = 8'h8d; ram[16'h2449] = 8'h06; ram[16'h244a] = 8'h02; ram[16'h244b] = 8'h38; ram[16'h244c] = 8'h20; ram[16'h244d] = 8'hf7; ram[16'h244e] = 8'h24; ram[16'h244f] = 8'hc6; 
ram[16'h2450] = 8'h0c; ram[16'h2451] = 8'ha5; ram[16'h2452] = 8'h0f; ram[16'h2453] = 8'hd0; ram[16'h2454] = 8'h08; ram[16'h2455] = 8'hc6; ram[16'h2456] = 8'h10; ram[16'h2457] = 8'ha9; 
ram[16'h2458] = 8'h99; ram[16'h2459] = 8'h85; ram[16'h245a] = 8'h0f; ram[16'h245b] = 8'hd0; ram[16'h245c] = 8'h12; ram[16'h245d] = 8'h29; ram[16'h245e] = 8'h0f; ram[16'h245f] = 8'hd0; 

ram[16'h2460] = 8'h0c; ram[16'h2461] = 8'hc6; ram[16'h2462] = 8'h0f; ram[16'h2463] = 8'hc6; ram[16'h2464] = 8'h0f; ram[16'h2465] = 8'hc6; ram[16'h2466] = 8'h0f; ram[16'h2467] = 8'hc6; 
ram[16'h2468] = 8'h0f; ram[16'h2469] = 8'hc6; ram[16'h246a] = 8'h0f; ram[16'h246b] = 8'hc6; ram[16'h246c] = 8'h0f; ram[16'h246d] = 8'hc6; ram[16'h246e] = 8'h0f; ram[16'h246f] = 8'h08; 
ram[16'h2470] = 8'h68; ram[16'h2471] = 8'h29; ram[16'h2472] = 8'h82; ram[16'h2473] = 8'h05; ram[16'h2474] = 8'h10; ram[16'h2475] = 8'h85; ram[16'h2476] = 8'h11; ram[16'h2477] = 8'h18; 
ram[16'h2478] = 8'h20; ram[16'h2479] = 8'hf7; ram[16'h247a] = 8'h24; ram[16'h247b] = 8'he6; ram[16'h247c] = 8'h0c; ram[16'h247d] = 8'ha5; ram[16'h247e] = 8'h0d; ram[16'h247f] = 8'hf0; 

ram[16'h2480] = 8'h15; ram[16'h2481] = 8'h29; ram[16'h2482] = 8'h0f; ram[16'h2483] = 8'hd0; ram[16'h2484] = 8'h0c; ram[16'h2485] = 8'hc6; ram[16'h2486] = 8'h0d; ram[16'h2487] = 8'hc6; 
ram[16'h2488] = 8'h0d; ram[16'h2489] = 8'hc6; ram[16'h248a] = 8'h0d; ram[16'h248b] = 8'hc6; ram[16'h248c] = 8'h0d; ram[16'h248d] = 8'hc6; ram[16'h248e] = 8'h0d; ram[16'h248f] = 8'hc6; 
ram[16'h2490] = 8'h0d; ram[16'h2491] = 8'hc6; ram[16'h2492] = 8'h0d; ram[16'h2493] = 8'h4c; ram[16'h2494] = 8'h4b; ram[16'h2495] = 8'h24; ram[16'h2496] = 8'ha9; ram[16'h2497] = 8'h99; 
ram[16'h2498] = 8'h85; ram[16'h2499] = 8'h0d; ram[16'h249a] = 8'ha5; ram[16'h249b] = 8'h0e; ram[16'h249c] = 8'hf0; ram[16'h249d] = 8'h39; ram[16'h249e] = 8'h29; ram[16'h249f] = 8'h0f; 

ram[16'h24a0] = 8'hd0; ram[16'h24a1] = 8'h18; ram[16'h24a2] = 8'hc6; ram[16'h24a3] = 8'h0e; ram[16'h24a4] = 8'hc6; ram[16'h24a5] = 8'h0e; ram[16'h24a6] = 8'hc6; ram[16'h24a7] = 8'h0e; 
ram[16'h24a8] = 8'hc6; ram[16'h24a9] = 8'h0e; ram[16'h24aa] = 8'hc6; ram[16'h24ab] = 8'h0e; ram[16'h24ac] = 8'hc6; ram[16'h24ad] = 8'h0e; ram[16'h24ae] = 8'he6; ram[16'h24af] = 8'h12; 
ram[16'h24b0] = 8'he6; ram[16'h24b1] = 8'h12; ram[16'h24b2] = 8'he6; ram[16'h24b3] = 8'h12; ram[16'h24b4] = 8'he6; ram[16'h24b5] = 8'h12; ram[16'h24b6] = 8'he6; ram[16'h24b7] = 8'h12; 
ram[16'h24b8] = 8'he6; ram[16'h24b9] = 8'h12; ram[16'h24ba] = 8'hc6; ram[16'h24bb] = 8'h0e; ram[16'h24bc] = 8'he6; ram[16'h24bd] = 8'h12; ram[16'h24be] = 8'ha5; ram[16'h24bf] = 8'h12; 

ram[16'h24c0] = 8'h8d; ram[16'h24c1] = 8'h06; ram[16'h24c2] = 8'h02; ram[16'h24c3] = 8'ha5; ram[16'h24c4] = 8'h0e; ram[16'h24c5] = 8'h8d; ram[16'h24c6] = 8'h05; ram[16'h24c7] = 8'h02; 
ram[16'h24c8] = 8'h85; ram[16'h24c9] = 8'h0f; ram[16'h24ca] = 8'h08; ram[16'h24cb] = 8'h68; ram[16'h24cc] = 8'h29; ram[16'h24cd] = 8'h82; ram[16'h24ce] = 8'h09; ram[16'h24cf] = 8'h01; 
ram[16'h24d0] = 8'h85; ram[16'h24d1] = 8'h11; ram[16'h24d2] = 8'he6; ram[16'h24d3] = 8'h10; ram[16'h24d4] = 8'h4c; ram[16'h24d5] = 8'h4b; ram[16'h24d6] = 8'h24; ram[16'h24d7] = 8'he0; 
ram[16'h24d8] = 8'h0e; ram[16'h24d9] = 8'hd0; ram[16'h24da] = 8'hfe; ram[16'h24db] = 8'hc0; ram[16'h24dc] = 8'hff; ram[16'h24dd] = 8'hd0; ram[16'h24de] = 8'hfe; ram[16'h24df] = 8'hba; 

ram[16'h24e0] = 8'he0; ram[16'h24e1] = 8'hff; ram[16'h24e2] = 8'hd0; ram[16'h24e3] = 8'hfe; ram[16'h24e4] = 8'hd8; ram[16'h24e5] = 8'had; ram[16'h24e6] = 8'h02; ram[16'h24e7] = 8'h02; 
ram[16'h24e8] = 8'hc9; ram[16'h24e9] = 8'h15; ram[16'h24ea] = 8'hd0; ram[16'h24eb] = 8'hfe; ram[16'h24ec] = 8'ha9; ram[16'h24ed] = 8'hf0; ram[16'h24ee] = 8'h8d; ram[16'h24ef] = 8'h02; 
ram[16'h24f0] = 8'h02; ram[16'h24f1] = 8'h4c; ram[16'h24f2] = 8'hf1; ram[16'h24f3] = 8'h24; ram[16'h24f4] = 8'h4c; ram[16'h24f5] = 8'h00; ram[16'h24f6] = 8'h04; ram[16'h24f7] = 8'h08; 
ram[16'h24f8] = 8'ha5; ram[16'h24f9] = 8'h0d; ram[16'h24fa] = 8'h65; ram[16'h24fb] = 8'h0e; ram[16'h24fc] = 8'h08; ram[16'h24fd] = 8'hc5; ram[16'h24fe] = 8'h0f; ram[16'h24ff] = 8'hd0; 

ram[16'h2500] = 8'hfe; ram[16'h2501] = 8'h68; ram[16'h2502] = 8'h29; ram[16'h2503] = 8'h83; ram[16'h2504] = 8'hc5; ram[16'h2505] = 8'h11; ram[16'h2506] = 8'hd0; ram[16'h2507] = 8'hfe; 
ram[16'h2508] = 8'h28; ram[16'h2509] = 8'h08; ram[16'h250a] = 8'ha5; ram[16'h250b] = 8'h0d; ram[16'h250c] = 8'he5; ram[16'h250d] = 8'h12; ram[16'h250e] = 8'h08; ram[16'h250f] = 8'hc5; 
ram[16'h2510] = 8'h0f; ram[16'h2511] = 8'hd0; ram[16'h2512] = 8'hfe; ram[16'h2513] = 8'h68; ram[16'h2514] = 8'h29; ram[16'h2515] = 8'h83; ram[16'h2516] = 8'hc5; ram[16'h2517] = 8'h11; 
ram[16'h2518] = 8'hd0; ram[16'h2519] = 8'hfe; ram[16'h251a] = 8'h28; ram[16'h251b] = 8'h08; ram[16'h251c] = 8'ha5; ram[16'h251d] = 8'h0d; ram[16'h251e] = 8'h6d; ram[16'h251f] = 8'h05; 

ram[16'h2520] = 8'h02; ram[16'h2521] = 8'h08; ram[16'h2522] = 8'hc5; ram[16'h2523] = 8'h0f; ram[16'h2524] = 8'hd0; ram[16'h2525] = 8'hfe; ram[16'h2526] = 8'h68; ram[16'h2527] = 8'h29; 
ram[16'h2528] = 8'h83; ram[16'h2529] = 8'hc5; ram[16'h252a] = 8'h11; ram[16'h252b] = 8'hd0; ram[16'h252c] = 8'hfe; ram[16'h252d] = 8'h28; ram[16'h252e] = 8'h08; ram[16'h252f] = 8'ha5; 
ram[16'h2530] = 8'h0d; ram[16'h2531] = 8'hed; ram[16'h2532] = 8'h06; ram[16'h2533] = 8'h02; ram[16'h2534] = 8'h08; ram[16'h2535] = 8'hc5; ram[16'h2536] = 8'h0f; ram[16'h2537] = 8'hd0; 
ram[16'h2538] = 8'hfe; ram[16'h2539] = 8'h68; ram[16'h253a] = 8'h29; ram[16'h253b] = 8'h83; ram[16'h253c] = 8'hc5; ram[16'h253d] = 8'h11; ram[16'h253e] = 8'hd0; ram[16'h253f] = 8'hfe; 

ram[16'h2540] = 8'h28; ram[16'h2541] = 8'h08; ram[16'h2542] = 8'ha5; ram[16'h2543] = 8'h0e; ram[16'h2544] = 8'h8d; ram[16'h2545] = 8'h0b; ram[16'h2546] = 8'h02; ram[16'h2547] = 8'ha5; 
ram[16'h2548] = 8'h0d; ram[16'h2549] = 8'h20; ram[16'h254a] = 8'h0a; ram[16'h254b] = 8'h02; ram[16'h254c] = 8'h08; ram[16'h254d] = 8'hc5; ram[16'h254e] = 8'h0f; ram[16'h254f] = 8'hd0; 
ram[16'h2550] = 8'hfe; ram[16'h2551] = 8'h68; ram[16'h2552] = 8'h29; ram[16'h2553] = 8'h83; ram[16'h2554] = 8'hc5; ram[16'h2555] = 8'h11; ram[16'h2556] = 8'hd0; ram[16'h2557] = 8'hfe; 
ram[16'h2558] = 8'h28; ram[16'h2559] = 8'h08; ram[16'h255a] = 8'ha5; ram[16'h255b] = 8'h12; ram[16'h255c] = 8'h8d; ram[16'h255d] = 8'h0e; ram[16'h255e] = 8'h02; ram[16'h255f] = 8'ha5; 

ram[16'h2560] = 8'h0d; ram[16'h2561] = 8'h20; ram[16'h2562] = 8'h0d; ram[16'h2563] = 8'h02; ram[16'h2564] = 8'h08; ram[16'h2565] = 8'hc5; ram[16'h2566] = 8'h0f; ram[16'h2567] = 8'hd0; 
ram[16'h2568] = 8'hfe; ram[16'h2569] = 8'h68; ram[16'h256a] = 8'h29; ram[16'h256b] = 8'h83; ram[16'h256c] = 8'hc5; ram[16'h256d] = 8'h11; ram[16'h256e] = 8'hd0; ram[16'h256f] = 8'hfe; 
ram[16'h2570] = 8'h28; ram[16'h2571] = 8'h08; ram[16'h2572] = 8'ha5; ram[16'h2573] = 8'h0d; ram[16'h2574] = 8'h75; ram[16'h2575] = 8'h00; ram[16'h2576] = 8'h08; ram[16'h2577] = 8'hc5; 
ram[16'h2578] = 8'h0f; ram[16'h2579] = 8'hd0; ram[16'h257a] = 8'hfe; ram[16'h257b] = 8'h68; ram[16'h257c] = 8'h29; ram[16'h257d] = 8'h83; ram[16'h257e] = 8'hc5; ram[16'h257f] = 8'h11; 

ram[16'h2580] = 8'hd0; ram[16'h2581] = 8'hfe; ram[16'h2582] = 8'h28; ram[16'h2583] = 8'h08; ram[16'h2584] = 8'ha5; ram[16'h2585] = 8'h0d; ram[16'h2586] = 8'hf5; ram[16'h2587] = 8'h04; 
ram[16'h2588] = 8'h08; ram[16'h2589] = 8'hc5; ram[16'h258a] = 8'h0f; ram[16'h258b] = 8'hd0; ram[16'h258c] = 8'hfe; ram[16'h258d] = 8'h68; ram[16'h258e] = 8'h29; ram[16'h258f] = 8'h83; 
ram[16'h2590] = 8'hc5; ram[16'h2591] = 8'h11; ram[16'h2592] = 8'hd0; ram[16'h2593] = 8'hfe; ram[16'h2594] = 8'h28; ram[16'h2595] = 8'h08; ram[16'h2596] = 8'ha5; ram[16'h2597] = 8'h0d; 
ram[16'h2598] = 8'h7d; ram[16'h2599] = 8'hf7; ram[16'h259a] = 8'h01; ram[16'h259b] = 8'h08; ram[16'h259c] = 8'hc5; ram[16'h259d] = 8'h0f; ram[16'h259e] = 8'hd0; ram[16'h259f] = 8'hfe; 

ram[16'h25a0] = 8'h68; ram[16'h25a1] = 8'h29; ram[16'h25a2] = 8'h83; ram[16'h25a3] = 8'hc5; ram[16'h25a4] = 8'h11; ram[16'h25a5] = 8'hd0; ram[16'h25a6] = 8'hfe; ram[16'h25a7] = 8'h28; 
ram[16'h25a8] = 8'h08; ram[16'h25a9] = 8'ha5; ram[16'h25aa] = 8'h0d; ram[16'h25ab] = 8'hfd; ram[16'h25ac] = 8'hf8; ram[16'h25ad] = 8'h01; ram[16'h25ae] = 8'h08; ram[16'h25af] = 8'hc5; 
ram[16'h25b0] = 8'h0f; ram[16'h25b1] = 8'hd0; ram[16'h25b2] = 8'hfe; ram[16'h25b3] = 8'h68; ram[16'h25b4] = 8'h29; ram[16'h25b5] = 8'h83; ram[16'h25b6] = 8'hc5; ram[16'h25b7] = 8'h11; 
ram[16'h25b8] = 8'hd0; ram[16'h25b9] = 8'hfe; ram[16'h25ba] = 8'h28; ram[16'h25bb] = 8'h08; ram[16'h25bc] = 8'ha5; ram[16'h25bd] = 8'h0d; ram[16'h25be] = 8'h79; ram[16'h25bf] = 8'h06; 

ram[16'h25c0] = 8'h01; ram[16'h25c1] = 8'h08; ram[16'h25c2] = 8'hc5; ram[16'h25c3] = 8'h0f; ram[16'h25c4] = 8'hd0; ram[16'h25c5] = 8'hfe; ram[16'h25c6] = 8'h68; ram[16'h25c7] = 8'h29; 
ram[16'h25c8] = 8'h83; ram[16'h25c9] = 8'hc5; ram[16'h25ca] = 8'h11; ram[16'h25cb] = 8'hd0; ram[16'h25cc] = 8'hfe; ram[16'h25cd] = 8'h28; ram[16'h25ce] = 8'h08; ram[16'h25cf] = 8'ha5; 
ram[16'h25d0] = 8'h0d; ram[16'h25d1] = 8'hf9; ram[16'h25d2] = 8'h07; ram[16'h25d3] = 8'h01; ram[16'h25d4] = 8'h08; ram[16'h25d5] = 8'hc5; ram[16'h25d6] = 8'h0f; ram[16'h25d7] = 8'hd0; 
ram[16'h25d8] = 8'hfe; ram[16'h25d9] = 8'h68; ram[16'h25da] = 8'h29; ram[16'h25db] = 8'h83; ram[16'h25dc] = 8'hc5; ram[16'h25dd] = 8'h11; ram[16'h25de] = 8'hd0; ram[16'h25df] = 8'hfe; 

ram[16'h25e0] = 8'h28; ram[16'h25e1] = 8'h08; ram[16'h25e2] = 8'ha5; ram[16'h25e3] = 8'h0d; ram[16'h25e4] = 8'h61; ram[16'h25e5] = 8'h44; ram[16'h25e6] = 8'h08; ram[16'h25e7] = 8'hc5; 
ram[16'h25e8] = 8'h0f; ram[16'h25e9] = 8'hd0; ram[16'h25ea] = 8'hfe; ram[16'h25eb] = 8'h68; ram[16'h25ec] = 8'h29; ram[16'h25ed] = 8'h83; ram[16'h25ee] = 8'hc5; ram[16'h25ef] = 8'h11; 
ram[16'h25f0] = 8'hd0; ram[16'h25f1] = 8'hfe; ram[16'h25f2] = 8'h28; ram[16'h25f3] = 8'h08; ram[16'h25f4] = 8'ha5; ram[16'h25f5] = 8'h0d; ram[16'h25f6] = 8'he1; ram[16'h25f7] = 8'h46; 
ram[16'h25f8] = 8'h08; ram[16'h25f9] = 8'hc5; ram[16'h25fa] = 8'h0f; ram[16'h25fb] = 8'hd0; ram[16'h25fc] = 8'hfe; ram[16'h25fd] = 8'h68; ram[16'h25fe] = 8'h29; ram[16'h25ff] = 8'h83; 

ram[16'h2600] = 8'hc5; ram[16'h2601] = 8'h11; ram[16'h2602] = 8'hd0; ram[16'h2603] = 8'hfe; ram[16'h2604] = 8'h28; ram[16'h2605] = 8'h08; ram[16'h2606] = 8'ha5; ram[16'h2607] = 8'h0d; 
ram[16'h2608] = 8'h71; ram[16'h2609] = 8'h56; ram[16'h260a] = 8'h08; ram[16'h260b] = 8'hc5; ram[16'h260c] = 8'h0f; ram[16'h260d] = 8'hd0; ram[16'h260e] = 8'hfe; ram[16'h260f] = 8'h68; 
ram[16'h2610] = 8'h29; ram[16'h2611] = 8'h83; ram[16'h2612] = 8'hc5; ram[16'h2613] = 8'h11; ram[16'h2614] = 8'hd0; ram[16'h2615] = 8'hfe; ram[16'h2616] = 8'h28; ram[16'h2617] = 8'h08; 
ram[16'h2618] = 8'ha5; ram[16'h2619] = 8'h0d; ram[16'h261a] = 8'hf1; ram[16'h261b] = 8'h58; ram[16'h261c] = 8'h08; ram[16'h261d] = 8'hc5; ram[16'h261e] = 8'h0f; ram[16'h261f] = 8'hd0; 

ram[16'h2620] = 8'hfe; ram[16'h2621] = 8'h68; ram[16'h2622] = 8'h29; ram[16'h2623] = 8'h83; ram[16'h2624] = 8'hc5; ram[16'h2625] = 8'h11; ram[16'h2626] = 8'hd0; ram[16'h2627] = 8'hfe; 
ram[16'h2628] = 8'h28; ram[16'h2629] = 8'h08; ram[16'h262a] = 8'ha5; ram[16'h262b] = 8'h0d; ram[16'h262c] = 8'h72; ram[16'h262d] = 8'h52; ram[16'h262e] = 8'h08; ram[16'h262f] = 8'hc5; 
ram[16'h2630] = 8'h0f; ram[16'h2631] = 8'hd0; ram[16'h2632] = 8'hfe; ram[16'h2633] = 8'h68; ram[16'h2634] = 8'h29; ram[16'h2635] = 8'h83; ram[16'h2636] = 8'hc5; ram[16'h2637] = 8'h11; 
ram[16'h2638] = 8'hd0; ram[16'h2639] = 8'hfe; ram[16'h263a] = 8'h28; ram[16'h263b] = 8'h08; ram[16'h263c] = 8'ha5; ram[16'h263d] = 8'h0d; ram[16'h263e] = 8'hf2; ram[16'h263f] = 8'h54; 

ram[16'h2640] = 8'h08; ram[16'h2641] = 8'hc5; ram[16'h2642] = 8'h0f; ram[16'h2643] = 8'hd0; ram[16'h2644] = 8'hfe; ram[16'h2645] = 8'h68; ram[16'h2646] = 8'h29; ram[16'h2647] = 8'h83; 
ram[16'h2648] = 8'hc5; ram[16'h2649] = 8'h11; ram[16'h264a] = 8'hd0; ram[16'h264b] = 8'hfe; ram[16'h264c] = 8'h28; ram[16'h264d] = 8'h60; ram[16'h264e] = 8'ha5; ram[16'h264f] = 8'h11; 
ram[16'h2650] = 8'h29; ram[16'h2651] = 8'h83; ram[16'h2652] = 8'h48; ram[16'h2653] = 8'ha5; ram[16'h2654] = 8'h0d; ram[16'h2655] = 8'h45; ram[16'h2656] = 8'h0e; ram[16'h2657] = 8'h30; 
ram[16'h2658] = 8'h0a; ram[16'h2659] = 8'ha5; ram[16'h265a] = 8'h0d; ram[16'h265b] = 8'h45; ram[16'h265c] = 8'h0f; ram[16'h265d] = 8'h10; ram[16'h265e] = 8'h04; ram[16'h265f] = 8'h68; 

ram[16'h2660] = 8'h09; ram[16'h2661] = 8'h40; ram[16'h2662] = 8'h48; ram[16'h2663] = 8'h68; ram[16'h2664] = 8'h85; ram[16'h2665] = 8'h11; ram[16'h2666] = 8'h08; ram[16'h2667] = 8'ha5; 
ram[16'h2668] = 8'h0d; ram[16'h2669] = 8'h72; ram[16'h266a] = 8'h52; ram[16'h266b] = 8'h08; ram[16'h266c] = 8'hc5; ram[16'h266d] = 8'h0f; ram[16'h266e] = 8'hd0; ram[16'h266f] = 8'hfe; 
ram[16'h2670] = 8'h68; ram[16'h2671] = 8'h29; ram[16'h2672] = 8'hc3; ram[16'h2673] = 8'hc5; ram[16'h2674] = 8'h11; ram[16'h2675] = 8'hd0; ram[16'h2676] = 8'hfe; ram[16'h2677] = 8'h28; 
ram[16'h2678] = 8'h08; ram[16'h2679] = 8'ha5; ram[16'h267a] = 8'h0d; ram[16'h267b] = 8'hf2; ram[16'h267c] = 8'h54; ram[16'h267d] = 8'h08; ram[16'h267e] = 8'hc5; ram[16'h267f] = 8'h0f; 

ram[16'h2680] = 8'hd0; ram[16'h2681] = 8'hfe; ram[16'h2682] = 8'h68; ram[16'h2683] = 8'h29; ram[16'h2684] = 8'hc3; ram[16'h2685] = 8'hc5; ram[16'h2686] = 8'h11; ram[16'h2687] = 8'hd0; 
ram[16'h2688] = 8'hfe; ram[16'h2689] = 8'h28; ram[16'h268a] = 8'h60; ram[16'h268b] = 8'h91; ram[16'h268c] = 8'h26; ram[16'h268d] = 8'h82; ram[16'h268e] = 8'h16; ram[16'h268f] = 8'h88; 
ram[16'h2690] = 8'h88; ram[16'h2691] = 8'h08; ram[16'h2692] = 8'h88; ram[16'h2693] = 8'h88; ram[16'h2694] = 8'h88; ram[16'h2695] = 8'h28; ram[16'h2696] = 8'hb0; ram[16'h2697] = 8'hfe; 
ram[16'h2698] = 8'h70; ram[16'h2699] = 8'hfe; ram[16'h269a] = 8'h30; ram[16'h269b] = 8'hfe; ram[16'h269c] = 8'hf0; ram[16'h269d] = 8'hfe; ram[16'h269e] = 8'hc9; ram[16'h269f] = 8'h49; 

ram[16'h26a0] = 8'hd0; ram[16'h26a1] = 8'hfe; ram[16'h26a2] = 8'he0; ram[16'h26a3] = 8'h4e; ram[16'h26a4] = 8'hd0; ram[16'h26a5] = 8'hfe; ram[16'h26a6] = 8'hc0; ram[16'h26a7] = 8'h41; 
ram[16'h26a8] = 8'hd0; ram[16'h26a9] = 8'hfe; ram[16'h26aa] = 8'h48; ram[16'h26ab] = 8'h8a; ram[16'h26ac] = 8'h48; ram[16'h26ad] = 8'hba; ram[16'h26ae] = 8'he0; ram[16'h26af] = 8'hfd; 
ram[16'h26b0] = 8'hd0; ram[16'h26b1] = 8'hfe; ram[16'h26b2] = 8'h68; ram[16'h26b3] = 8'haa; ram[16'h26b4] = 8'ha9; ram[16'h26b5] = 8'hff; ram[16'h26b6] = 8'h48; ram[16'h26b7] = 8'h28; 
ram[16'h26b8] = 8'h68; ram[16'h26b9] = 8'he8; ram[16'h26ba] = 8'h49; ram[16'h26bb] = 8'haa; ram[16'h26bc] = 8'h6c; ram[16'h26bd] = 8'hff; ram[16'h26be] = 8'h02; ram[16'h26bf] = 8'hea; 

ram[16'h26c0] = 8'hea; ram[16'h26c1] = 8'h4c; ram[16'h26c2] = 8'hc1; ram[16'h26c3] = 8'h26; ram[16'h26c4] = 8'h4c; ram[16'h26c5] = 8'h00; ram[16'h26c6] = 8'h04; ram[16'h26c7] = 8'h0e; 
ram[16'h26c8] = 8'h27; ram[16'h26c9] = 8'h0e; ram[16'h26ca] = 8'h27; ram[16'h26cb] = 8'hd5; ram[16'h26cc] = 8'h26; ram[16'h26cd] = 8'hce; ram[16'h26ce] = 8'h16; ram[16'h26cf] = 8'h0e; 
ram[16'h26d0] = 8'h27; ram[16'h26d1] = 8'h0e; ram[16'h26d2] = 8'h27; ram[16'h26d3] = 8'h88; ram[16'h26d4] = 8'h88; ram[16'h26d5] = 8'h08; ram[16'h26d6] = 8'h88; ram[16'h26d7] = 8'h88; 
ram[16'h26d8] = 8'h88; ram[16'h26d9] = 8'h28; ram[16'h26da] = 8'hb0; ram[16'h26db] = 8'hfe; ram[16'h26dc] = 8'h70; ram[16'h26dd] = 8'hfe; ram[16'h26de] = 8'h30; ram[16'h26df] = 8'hfe; 

ram[16'h26e0] = 8'hf0; ram[16'h26e1] = 8'hfe; ram[16'h26e2] = 8'hc9; ram[16'h26e3] = 8'h58; ram[16'h26e4] = 8'hd0; ram[16'h26e5] = 8'hfe; ram[16'h26e6] = 8'he0; ram[16'h26e7] = 8'h04; 
ram[16'h26e8] = 8'hd0; ram[16'h26e9] = 8'hfe; ram[16'h26ea] = 8'hc0; ram[16'h26eb] = 8'h46; ram[16'h26ec] = 8'hd0; ram[16'h26ed] = 8'hfe; ram[16'h26ee] = 8'h48; ram[16'h26ef] = 8'h8a; 
ram[16'h26f0] = 8'h48; ram[16'h26f1] = 8'hba; ram[16'h26f2] = 8'he0; ram[16'h26f3] = 8'hfd; ram[16'h26f4] = 8'hd0; ram[16'h26f5] = 8'hfe; ram[16'h26f6] = 8'h68; ram[16'h26f7] = 8'haa; 
ram[16'h26f8] = 8'ha9; ram[16'h26f9] = 8'hff; ram[16'h26fa] = 8'h48; ram[16'h26fb] = 8'h28; ram[16'h26fc] = 8'h68; ram[16'h26fd] = 8'he8; ram[16'h26fe] = 8'he8; ram[16'h26ff] = 8'h49; 

ram[16'h2700] = 8'haa; ram[16'h2701] = 8'h7c; ram[16'h2702] = 8'hf9; ram[16'h2703] = 8'h02; ram[16'h2704] = 8'hea; ram[16'h2705] = 8'hea; ram[16'h2706] = 8'h4c; ram[16'h2707] = 8'h06; 
ram[16'h2708] = 8'h27; ram[16'h2709] = 8'h4c; ram[16'h270a] = 8'h00; ram[16'h270b] = 8'h04; ram[16'h270c] = 8'hea; ram[16'h270d] = 8'hea; ram[16'h270e] = 8'hea; ram[16'h270f] = 8'hea; 
ram[16'h2710] = 8'h4c; ram[16'h2711] = 8'h10; ram[16'h2712] = 8'h27; ram[16'h2713] = 8'h4c; ram[16'h2714] = 8'h00; ram[16'h2715] = 8'h04; ram[16'h2716] = 8'h4c; ram[16'h2717] = 8'h16; 
ram[16'h2718] = 8'h27; ram[16'h2719] = 8'h4c; ram[16'h271a] = 8'h00; ram[16'h271b] = 8'h04; ram[16'h271c] = 8'h4c; ram[16'h271d] = 8'h1c; ram[16'h271e] = 8'h27; ram[16'h271f] = 8'h4c; 

ram[16'h2720] = 8'h00; ram[16'h2721] = 8'h04; ram[16'h2722] = 8'h88; ram[16'h2723] = 8'h88; ram[16'h2724] = 8'h08; ram[16'h2725] = 8'h88; ram[16'h2726] = 8'h88; ram[16'h2727] = 8'h88; 
ram[16'h2728] = 8'hc9; ram[16'h2729] = 8'hbd; ram[16'h272a] = 8'hf0; ram[16'h272b] = 8'h42; ram[16'h272c] = 8'hc9; ram[16'h272d] = 8'h42; ram[16'h272e] = 8'hd0; ram[16'h272f] = 8'hfe; 
ram[16'h2730] = 8'he0; ram[16'h2731] = 8'h52; ram[16'h2732] = 8'hd0; ram[16'h2733] = 8'hfe; ram[16'h2734] = 8'hc0; ram[16'h2735] = 8'h48; ram[16'h2736] = 8'hd0; ram[16'h2737] = 8'hfe; 
ram[16'h2738] = 8'h85; ram[16'h2739] = 8'h0a; ram[16'h273a] = 8'h86; ram[16'h273b] = 8'h0b; ram[16'h273c] = 8'hba; ram[16'h273d] = 8'hbd; ram[16'h273e] = 8'h02; ram[16'h273f] = 8'h01; 

ram[16'h2740] = 8'hc9; ram[16'h2741] = 8'h30; ram[16'h2742] = 8'hd0; ram[16'h2743] = 8'hfe; ram[16'h2744] = 8'h68; ram[16'h2745] = 8'hc9; ram[16'h2746] = 8'h34; ram[16'h2747] = 8'hd0; 
ram[16'h2748] = 8'hfe; ram[16'h2749] = 8'hba; ram[16'h274a] = 8'he0; ram[16'h274b] = 8'hfc; ram[16'h274c] = 8'hd0; ram[16'h274d] = 8'hfe; ram[16'h274e] = 8'had; ram[16'h274f] = 8'hff; 
ram[16'h2750] = 8'h01; ram[16'h2751] = 8'hc9; ram[16'h2752] = 8'h17; ram[16'h2753] = 8'hd0; ram[16'h2754] = 8'hfe; ram[16'h2755] = 8'had; ram[16'h2756] = 8'hfe; ram[16'h2757] = 8'h01; 
ram[16'h2758] = 8'hc9; ram[16'h2759] = 8'h20; ram[16'h275a] = 8'hd0; ram[16'h275b] = 8'hfe; ram[16'h275c] = 8'ha9; ram[16'h275d] = 8'hff; ram[16'h275e] = 8'h48; ram[16'h275f] = 8'ha6; 

ram[16'h2760] = 8'h0b; ram[16'h2761] = 8'he8; ram[16'h2762] = 8'ha5; ram[16'h2763] = 8'h0a; ram[16'h2764] = 8'h49; ram[16'h2765] = 8'haa; ram[16'h2766] = 8'h28; ram[16'h2767] = 8'h40; 
ram[16'h2768] = 8'h4c; ram[16'h2769] = 8'h68; ram[16'h276a] = 8'h27; ram[16'h276b] = 8'h4c; ram[16'h276c] = 8'h00; ram[16'h276d] = 8'h04; ram[16'h276e] = 8'he0; ram[16'h276f] = 8'had; 
ram[16'h2770] = 8'hd0; ram[16'h2771] = 8'hfe; ram[16'h2772] = 8'hc0; ram[16'h2773] = 8'hb1; ram[16'h2774] = 8'hd0; ram[16'h2775] = 8'hfe; ram[16'h2776] = 8'h85; ram[16'h2777] = 8'h0a; 
ram[16'h2778] = 8'h86; ram[16'h2779] = 8'h0b; ram[16'h277a] = 8'hba; ram[16'h277b] = 8'hbd; ram[16'h277c] = 8'h02; ram[16'h277d] = 8'h01; ram[16'h277e] = 8'hc9; ram[16'h277f] = 8'hff; 

ram[16'h2780] = 8'hd0; ram[16'h2781] = 8'hfe; ram[16'h2782] = 8'h68; ram[16'h2783] = 8'hc9; ram[16'h2784] = 8'hf7; ram[16'h2785] = 8'hd0; ram[16'h2786] = 8'hfe; ram[16'h2787] = 8'hba; 
ram[16'h2788] = 8'he0; ram[16'h2789] = 8'hfc; ram[16'h278a] = 8'hd0; ram[16'h278b] = 8'hfe; ram[16'h278c] = 8'had; ram[16'h278d] = 8'hff; ram[16'h278e] = 8'h01; ram[16'h278f] = 8'hc9; 
ram[16'h2790] = 8'h17; ram[16'h2791] = 8'hd0; ram[16'h2792] = 8'hfe; ram[16'h2793] = 8'had; ram[16'h2794] = 8'hfe; ram[16'h2795] = 8'h01; ram[16'h2796] = 8'hc9; ram[16'h2797] = 8'h46; 
ram[16'h2798] = 8'hd0; ram[16'h2799] = 8'hfe; ram[16'h279a] = 8'ha9; ram[16'h279b] = 8'h04; ram[16'h279c] = 8'h48; ram[16'h279d] = 8'ha6; ram[16'h279e] = 8'h0b; ram[16'h279f] = 8'he8; 

ram[16'h27a0] = 8'ha5; ram[16'h27a1] = 8'h0a; ram[16'h27a2] = 8'h49; ram[16'h27a3] = 8'haa; ram[16'h27a4] = 8'h28; ram[16'h27a5] = 8'h40; ram[16'h27a6] = 8'h4c; ram[16'h27a7] = 8'ha6; 
ram[16'h27a8] = 8'h27; ram[16'h27a9] = 8'h4c; ram[16'h27aa] = 8'h00; ram[16'h27ab] = 8'h04; ram[16'h27ac] = 8'h00; ram[16'h27ad] = 8'h00; ram[16'h27ae] = 8'h00; ram[16'h27af] = 8'h00; 
ram[16'h27b0] = 8'h00; ram[16'h27b1] = 8'h00; ram[16'h27b2] = 8'h00; ram[16'h27b3] = 8'h00; ram[16'h27b4] = 8'h00; ram[16'h27b5] = 8'h00; ram[16'h27b6] = 8'h00; ram[16'h27b7] = 8'h00; 
ram[16'h27b8] = 8'h00; ram[16'h27b9] = 8'h00; ram[16'h27ba] = 8'h00; ram[16'h27bb] = 8'h00; ram[16'h27bc] = 8'h00; ram[16'h27bd] = 8'h00; ram[16'h27be] = 8'h00; ram[16'h27bf] = 8'h00; 

ram[16'h27c0] = 8'h00; ram[16'h27c1] = 8'h00; ram[16'h27c2] = 8'h00; ram[16'h27c3] = 8'h00; ram[16'h27c4] = 8'h00; ram[16'h27c5] = 8'h00; ram[16'h27c6] = 8'h00; ram[16'h27c7] = 8'h00; 
ram[16'h27c8] = 8'h00; ram[16'h27c9] = 8'h00; ram[16'h27ca] = 8'h00; ram[16'h27cb] = 8'h00; ram[16'h27cc] = 8'hea; ram[16'h27cd] = 8'hea; ram[16'h27ce] = 8'hea; ram[16'h27cf] = 8'hea; 
ram[16'h27d0] = 8'h4c; ram[16'h27d1] = 8'hd0; ram[16'h27d2] = 8'h27; ram[16'h27d3] = 8'h00; ram[16'h27d4] = 8'h00; ram[16'h27d5] = 8'h00; ram[16'h27d6] = 8'h00; ram[16'h27d7] = 8'h00; 
ram[16'h27d8] = 8'h00; ram[16'h27d9] = 8'h00; ram[16'h27da] = 8'h00; ram[16'h27db] = 8'h00; ram[16'h27dc] = 8'h00; ram[16'h27dd] = 8'h00; ram[16'h27de] = 8'h00; ram[16'h27df] = 8'h00; 

ram[16'h27e0] = 8'h00; ram[16'h27e1] = 8'h00; ram[16'h27e2] = 8'h00; ram[16'h27e3] = 8'h00; ram[16'h27e4] = 8'h00; ram[16'h27e5] = 8'h00; ram[16'h27e6] = 8'h00; ram[16'h27e7] = 8'h00; 
ram[16'h27e8] = 8'h00; ram[16'h27e9] = 8'h00; ram[16'h27ea] = 8'h00; ram[16'h27eb] = 8'h00; ram[16'h27ec] = 8'h00; ram[16'h27ed] = 8'h00; ram[16'h27ee] = 8'h00; ram[16'h27ef] = 8'h00; 
ram[16'h27f0] = 8'h00; ram[16'h27f1] = 8'h00; ram[16'h27f2] = 8'h00; ram[16'h27f3] = 8'h00; ram[16'h27f4] = 8'h00; ram[16'h27f5] = 8'h00; ram[16'h27f6] = 8'h00; ram[16'h27f7] = 8'h00; 
ram[16'h27f8] = 8'h00; ram[16'h27f9] = 8'h00; ram[16'h27fa] = 8'h00; ram[16'h27fb] = 8'h00; ram[16'h27fc] = 8'h00; ram[16'h27fd] = 8'h00; ram[16'h27fe] = 8'h00; ram[16'h27ff] = 8'h00; 

ram[16'h2800] = 8'h00; ram[16'h2801] = 8'h00; ram[16'h2802] = 8'h00; ram[16'h2803] = 8'h00; ram[16'h2804] = 8'h00; ram[16'h2805] = 8'h00; ram[16'h2806] = 8'h00; ram[16'h2807] = 8'h00; 
ram[16'h2808] = 8'h00; ram[16'h2809] = 8'h00; ram[16'h280a] = 8'h00; ram[16'h280b] = 8'h00; ram[16'h280c] = 8'h00; ram[16'h280d] = 8'h00; ram[16'h280e] = 8'h00; ram[16'h280f] = 8'h00; 
ram[16'h2810] = 8'h00; ram[16'h2811] = 8'h00; ram[16'h2812] = 8'h00; ram[16'h2813] = 8'h00; ram[16'h2814] = 8'h00; ram[16'h2815] = 8'h00; ram[16'h2816] = 8'h00; ram[16'h2817] = 8'h00; 
ram[16'h2818] = 8'h00; ram[16'h2819] = 8'h00; ram[16'h281a] = 8'h00; ram[16'h281b] = 8'h00; ram[16'h281c] = 8'h00; ram[16'h281d] = 8'h00; ram[16'h281e] = 8'h00; ram[16'h281f] = 8'h00; 

ram[16'h2820] = 8'h00; ram[16'h2821] = 8'h00; ram[16'h2822] = 8'h00; ram[16'h2823] = 8'h00; ram[16'h2824] = 8'h00; ram[16'h2825] = 8'h00; ram[16'h2826] = 8'h00; ram[16'h2827] = 8'h00; 
ram[16'h2828] = 8'h00; ram[16'h2829] = 8'h00; ram[16'h282a] = 8'h00; ram[16'h282b] = 8'h00; ram[16'h282c] = 8'h00; ram[16'h282d] = 8'h00; ram[16'h282e] = 8'h00; ram[16'h282f] = 8'h00; 
ram[16'h2830] = 8'h00; ram[16'h2831] = 8'h00; ram[16'h2832] = 8'h00; ram[16'h2833] = 8'h00; ram[16'h2834] = 8'h00; ram[16'h2835] = 8'h00; ram[16'h2836] = 8'h00; ram[16'h2837] = 8'h00; 
ram[16'h2838] = 8'h00; ram[16'h2839] = 8'h00; ram[16'h283a] = 8'h00; ram[16'h283b] = 8'h00; ram[16'h283c] = 8'h00; ram[16'h283d] = 8'h00; ram[16'h283e] = 8'h00; ram[16'h283f] = 8'h00; 

ram[16'h2840] = 8'h00; ram[16'h2841] = 8'h00; ram[16'h2842] = 8'h00; ram[16'h2843] = 8'h00; ram[16'h2844] = 8'h00; ram[16'h2845] = 8'h00; ram[16'h2846] = 8'h00; ram[16'h2847] = 8'h00; 
ram[16'h2848] = 8'h00; ram[16'h2849] = 8'h00; ram[16'h284a] = 8'h00; ram[16'h284b] = 8'h00; ram[16'h284c] = 8'h00; ram[16'h284d] = 8'h00; ram[16'h284e] = 8'h00; ram[16'h284f] = 8'h00; 
ram[16'h2850] = 8'h00; ram[16'h2851] = 8'h00; ram[16'h2852] = 8'h00; ram[16'h2853] = 8'h00; ram[16'h2854] = 8'h00; ram[16'h2855] = 8'h00; ram[16'h2856] = 8'h00; ram[16'h2857] = 8'h00; 
ram[16'h2858] = 8'h00; ram[16'h2859] = 8'h00; ram[16'h285a] = 8'h00; ram[16'h285b] = 8'h00; ram[16'h285c] = 8'h00; ram[16'h285d] = 8'h00; ram[16'h285e] = 8'h00; ram[16'h285f] = 8'h00; 

ram[16'h2860] = 8'h00; ram[16'h2861] = 8'h00; ram[16'h2862] = 8'h00; ram[16'h2863] = 8'h00; ram[16'h2864] = 8'h00; ram[16'h2865] = 8'h00; ram[16'h2866] = 8'h00; ram[16'h2867] = 8'h00; 
ram[16'h2868] = 8'h00; ram[16'h2869] = 8'h00; ram[16'h286a] = 8'h00; ram[16'h286b] = 8'h00; ram[16'h286c] = 8'h00; ram[16'h286d] = 8'h00; ram[16'h286e] = 8'h00; ram[16'h286f] = 8'h00; 
ram[16'h2870] = 8'h00; ram[16'h2871] = 8'h00; ram[16'h2872] = 8'h00; ram[16'h2873] = 8'h00; ram[16'h2874] = 8'h00; ram[16'h2875] = 8'h00; ram[16'h2876] = 8'h00; ram[16'h2877] = 8'h00; 
ram[16'h2878] = 8'h00; ram[16'h2879] = 8'h00; ram[16'h287a] = 8'h00; ram[16'h287b] = 8'h00; ram[16'h287c] = 8'h00; ram[16'h287d] = 8'h00; ram[16'h287e] = 8'h00; ram[16'h287f] = 8'h00; 

ram[16'h2880] = 8'hea; ram[16'h2881] = 8'hea; ram[16'h2882] = 8'hea; ram[16'h2883] = 8'hea; ram[16'h2884] = 8'h4c; ram[16'h2885] = 8'h84; ram[16'h2886] = 8'h28; 
ram[16'hfffa] = 8'h16; ram[16'hfffb] = 8'h27; ram[16'hfffc] = 8'h1c; ram[16'hfffd] = 8'h27; ram[16'hfffe] = 8'h24; ram[16'hffff] = 8'h27; 
 // Override start vector
ram[16'hfffc] = 8'h00;
ram[16'hfffd] = 8'h04;
end

always @(posedge clk)
begin
    if(we)
        ram[addr_w] = di;
    if(we && addr_w == 16'h0202)
        $display("last test: %d",di);
    do = ram[addr_r];
end

endmodule
